-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- 
-- ============================================================================
-- Module:					TODO
--
-- Authors:					Patrick Lehmann
-- 
-- Description:
-- ------------------------------------
--
-- Policies														| supported
-- -----------------------------------#--------------------
--	RR			round robin								| not yet
--	RAND		random										| not yet
--	CLOCK		clock algorithm						| not yet
--	LRU			least recently used				| YES
--	LFU			least frequently used			| not yet
-- -----------------------------------#--------------------
--
-- Priority		Command
-- ----------------------
--	0					invalidate
--	1					replace
--	2					access
--
-- License:
-- ============================================================================
-- Copyright 2007-2016 Technische Universitaet Dresden - Germany
--										 Chair for VLSI-Design, Diagnostics and Architecture
-- 
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
-- 
--		http://www.apache.org/licenses/LICENSE-2.0
-- 
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- ============================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

library PoC;
use PoC.config.all;
use PoC.utils.all;
use PoC.vectors.all;
use PoC.strings.all;


entity cache_replacement_policy is
	generic (
		REPLACEMENT_POLICY : string		:= "LRU";
		CACHE_LINES				 : positive := 32
	);
	port (
		Clock : in std_logic;
		Reset : in std_logic;

		-- replacement interface
		Replace			 : in	 std_logic;
		ReplaceIndex : out std_logic_vector(log2ceilnz(CACHE_LINES) - 1 downto 0);

		-- cacheline usage update interface
		TagAccess	 : in std_logic;
		ReadWrite	 : in std_logic;
		Invalidate : in std_logic;
		Index			 : in std_logic_vector(log2ceilnz(CACHE_LINES) - 1 downto 0)
	);
end;


architecture rtl of cache_replacement_policy is
	attribute KEEP				 : boolean;
	attribute FSM_ENCODING : string;

	constant KEY_BITS : positive := log2ceilnz(CACHE_LINES);

begin
	assert (str_equal(REPLACEMENT_POLICY, "RR") or
					str_equal(REPLACEMENT_POLICY, "LRU"))
		report "Unsupported replacement strategy"
		severity error;


	-- ===========================================================================
	-- policy: RR - round robin
	-- ===========================================================================
	genRR : if (str_equal(REPLACEMENT_POLICY, "RR") = true) generate
		constant VALID_BIT : natural := 0;

		subtype T_OPTION_LINE is std_logic_vector(0 downto 0);
		type T_OPTION_LINE_VECTOR is array (natural range <>) of T_OPTION_LINE;

		signal OptionMemory : T_OPTION_LINE_VECTOR(CACHE_LINES - 1 downto 0) := (others => (
			VALID_BIT																																			=> '0')
																																						 );

		signal ValidHit		: std_logic;
		signal Pointer_us : unsigned(log2ceilnz(CACHE_LINES) - 1 downto 0) := (others => '0');

	begin
--		ValidHit		<= OptionMemory(to_integer(unsigned(Index)))(VALID_BIT);
--		IsValid			<= ValidHit;
--
--		PROCESS(Clock)
--		BEGIN
--			IF rising_edge(Clock) THEN
--				IF (Reset = '1') THEN
--					FOR I IN 0 TO CACHE_LINES - 1 LOOP
--						OptionMemory(I)(VALID_BIT)	<= '0';
--					END LOOP;
--				ELSE
--					IF (Insert = '1') THEN
--						OptionMemory(to_integer(Pointer_us))(VALID_BIT) <= '1';
--					END IF;
--					
--					IF (Invalidate = '1') THEN
--						OptionMemory(to_integer(unsigned(Index)))(VALID_BIT)			<= '0';
--					END IF;
--				END IF;
--			END IF;
--		END PROCESS;
--
--		Replace				<= Insert;
--		ReplaceIndex	<= std_logic_vector(Pointer_us);
--		
--		PROCESS(Clock)
--		BEGIN
--			IF rising_edge(Clock) THEN
--				IF (Reset = '1') THEN
--					Pointer_us		<= (OTHERS => '0');
--				ELSE
--					IF (Insert = '1') THEN
--						Pointer_us	<= Pointer_us + 1;
--					END IF;
--				END IF;
--			END IF;
--		END PROCESS;
	end generate;

	-- ===========================================================================
	-- policy: LRU - least recently used
	-- ===========================================================================
	genLRU : if (str_equal(REPLACEMENT_POLICY, "LRU") = true) generate
		signal LRU_Insert			: std_logic;
		signal LRU_Invalidate : std_logic;
		signal KeyIn					: std_logic_vector(log2ceilnz(CACHE_LINES) - 1 downto 0);
		signal LRU_Key				: std_logic_vector(log2ceilnz(CACHE_LINES) - 1 downto 0);

	begin
		-- list_lru_systolic supports only one update per cycle
		process(TagAccess, ReadWrite, Invalidate, Replace, Index, LRU_Key)
		begin
			LRU_Insert		 <= '0';
			LRU_Invalidate <= '0';
			KeyIn					 <= Index;

			if (Invalidate = '1') then
				LRU_Invalidate <= '1';
				KeyIn					 <= Index;
			elsif (Replace = '1') then
				LRU_Insert <= '1';
				KeyIn			 <= LRU_Key;
			elsif (TagAccess = '1') then
				LRU_Insert <= '1';
				KeyIn			 <= Index;
			end if;
		end process;

		ReplaceIndex <= LRU_Key;

		LRU : entity PoC.sort_lru_cache
			generic map (
				ELEMENTS => CACHE_LINES
			)
			port map (
				Clock => Clock,
				Reset => Reset,

				Insert => LRU_Insert,
				Free	 => LRU_Invalidate,
				KeyIn	 => KeyIn,

				KeyOut => LRU_Key
			);
	end generate;
end architecture;
