-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- =============================================================================
-- Authors:					Patrick Lehmann
--									Martin Zabel
--
-- Entity:					OOB Sequencer for SATA Physical Layer - Device Side
--
-- Description:
-- -------------------------------------
-- Executes the COMRESET / COMINIT procedure.
--
-- If the clock is unstable, than Reset must be asserted.
-- Automatically tries to establish a communication when Reset is deasserted.
--
-- License:
-- =============================================================================
-- Copyright 2007-2015 Technische Universitaet Dresden - Germany
--										 Chair for VLSI-Design, Diagnostics and Architecture
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--		http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- =============================================================================

library IEEE;
use			IEEE.STD_LOGIC_1164.all;
use			IEEE.NUMERIC_STD.all;

library PoC;
use			PoC.config.all;
use			PoC.utils.all;
use			PoC.vectors.all;
use			PoC.strings.all;
use			PoC.physical.all;
use			PoC.debug.all;
use			PoC.sata.all;
use			PoC.satadbg.all;


entity sata_Physical_OOBControl_Device is
	generic (
		DEBUG											: boolean														:= FALSE;												-- generate additional debug signals and preserve them (attribute keep)
		ENABLE_DEBUGPORT					: boolean														:= FALSE;												-- enables the assignment of signals to the debugport
		ALLOW_STANDARD_VIOLATION	: boolean														:= FALSE;
		OOB_TIMEOUT								: T_TIME														:= T_TIME'low
	);
	port (
		Clock											: in	std_logic;
		Reset											: in	std_logic;
		-- debug ports
		DebugPortOut							: out	T_SATADBG_PHYSICAL_OOBCONTROL_OUT;

		Timeout										: out	std_logic;
		SATAGeneration						: in	T_SATA_GENERATION;
		HostDetected							: out	std_logic;
		LinkOK										: out	std_logic;
		LinkDead									: out	std_logic;

		OOB_TX_Command						: out	T_SATA_OOB;
		OOB_TX_Complete						: in	std_logic;
		OOB_RX_Received						: in	T_SATA_OOB;
		OOB_HandshakeComplete			:	out	std_logic;

		TX_Primitive							: out	T_SATA_PRIMITIVE;
		RX_Primitive							: in	T_SATA_PRIMITIVE;
		RX_Valid									: in	std_logic
	);
end entity;


architecture rtl of sata_Physical_OOBControl_Device is
	attribute KEEP												: boolean;
	attribute FSM_ENCODING								: string;

	constant CLOCK_GEN1_FREQ							: FREQ				:= 37500 kHz;		-- SATAClock frequency for SATA generation 1
	constant CLOCK_GEN2_FREQ							: FREQ				:= 75 MHz;			-- SATAClock frequency for SATA generation 2
	constant CLOCK_GEN3_FREQ							: FREQ				:= 150 MHz;			-- SATAClock frequency for SATA generation 3

	constant DEFAULT_OOB_TIMEOUT					: T_TIME			:= 880.0e-6;

	constant OOB_TIMEOUT_I								: T_TIME			:= ite((OOB_TIMEOUT = T_TIME'low), DEFAULT_OOB_TIMEOUT, OOB_TIMEOUT);
	constant COMRESET_TIMEOUT							: T_TIME			:= 450.0e-9;
	constant COMWAKE_TIMEOUT							: T_TIME			:= 250.0e-9;

	constant TTID1_OOB_TIMEOUT_GEN1				: natural			:= 0;
	constant TTID1_OOB_TIMEOUT_GEN2				: natural			:= 1;
	constant TTID1_OOB_TIMEOUT_GEN3				: natural			:= 2;
	constant TTID2_COMRESET_TIMEOUT_GEN1	: natural			:= 0;
	constant TTID2_COMRESET_TIMEOUT_GEN2	: natural			:= 1;
	constant TTID2_COMRESET_TIMEOUT_GEN3	: natural			:= 2;
	constant TTID2_COMWAKE_TIMEOUT_GEN1		: natural			:= 3;
	constant TTID2_COMWAKE_TIMEOUT_GEN2		: natural			:= 4;
	constant TTID2_COMWAKE_TIMEOUT_GEN3		: natural			:= 5;

	constant TC1_TIMING_TABLE					: T_NATVEC				:= (--		 880 us
		TTID1_OOB_TIMEOUT_GEN1 => TimingToCycles(OOB_TIMEOUT_I,	CLOCK_GEN1_FREQ),							-- slot 0
		TTID1_OOB_TIMEOUT_GEN2 => TimingToCycles(OOB_TIMEOUT_I,	CLOCK_GEN2_FREQ),							-- slot 1
		TTID1_OOB_TIMEOUT_GEN3 => TimingToCycles(OOB_TIMEOUT_I,	CLOCK_GEN3_FREQ)							-- slot 2
	);

	constant TC2_TIMING_TABLE					: T_NATVEC				:= (
		TTID2_COMRESET_TIMEOUT_GEN1	=> TimingToCycles(COMRESET_TIMEOUT,	CLOCK_GEN1_FREQ),		-- slot 0
		TTID2_COMRESET_TIMEOUT_GEN2	=> TimingToCycles(COMRESET_TIMEOUT,	CLOCK_GEN2_FREQ),		-- slot 1
		TTID2_COMRESET_TIMEOUT_GEN3	=> TimingToCycles(COMRESET_TIMEOUT,	CLOCK_GEN3_FREQ),		-- slot 2
		TTID2_COMWAKE_TIMEOUT_GEN1	=> TimingToCycles(COMWAKE_TIMEOUT,	CLOCK_GEN1_FREQ),		-- slot 3
		TTID2_COMWAKE_TIMEOUT_GEN2	=> TimingToCycles(COMWAKE_TIMEOUT,	CLOCK_GEN2_FREQ),		-- slot 4
		TTID2_COMWAKE_TIMEOUT_GEN3	=> TimingToCycles(COMWAKE_TIMEOUT,	CLOCK_GEN3_FREQ)		-- slot 5
	);

	type T_STATE is (
		ST_DEV_RESET,
		ST_DEV_WAIT_HOST_COMRESET,
		ST_DEV_WAIT_AFTER_HOST_COMRESET,
		ST_DEV_SEND_COMINIT,
		ST_DEV_WAIT_HOST_COMWAKE,
		ST_DEV_WAIT_AFTER_COMWAKE,
		ST_DEV_SEND_COMWAKE,
		ST_DEV_OOB_HANDSHAKE_COMPLETE,
		ST_DEV_SEND_ALIGN,
		ST_DEV_TIMEOUT,
		ST_DEV_LINK_OK,
		ST_DEV_LINK_DEAD
	);

	-- OOB-Statemachine
	signal State											: T_STATE														:= ST_DEV_RESET;
	signal NextState									: T_STATE;
	attribute FSM_ENCODING of State		: signal is getFSMEncoding_gray(DEBUG);

	signal HostDetected_i							: std_logic;
	signal LinkOK_i										: std_logic;
	signal LinkDead_i									: std_logic;
	signal Timeout_i									: std_logic;
	signal ReceivedReset_i						: std_logic;

	signal OOB_TX_Command_i						: T_SATA_OOB;
	signal OOB_HandshakeComplete_i		: std_logic;

	-- Timing-Counter
	-- ===========================================================================
	-- general timeouts
	signal TC1_en										: std_logic;
	signal TC1_Load									: std_logic;
	signal TC1_Slot									: natural;
	signal TC1_Timeout							: std_logic;

	-- OOB state specific timeouts
	signal TC2_en										: std_logic;
	signal TC2_Load									: std_logic;
	signal TC2_Slot									: natural;
	signal TC2_Timeout							: std_logic;

begin
	assert ((SATAGeneration = SATA_GENERATION_1) or
					(SATAGeneration = SATA_GENERATION_2) or
					(SATAGeneration = SATA_GENERATION_3))
		report "Member of T_SATA_GENERATION not supported"
		severity FAILURE;

	-- OOBControl Statemachine
	-- ======================================================================================================================================
	process(Clock)
	begin
		if rising_edge(Clock) then
			if (Reset = '1') then
				State			<= ST_DEV_RESET;
			else
				State			<= NextState;
			end if;
		end if;
	end process;


	process(State, SATAGeneration, OOB_TX_Complete, OOB_RX_Received, RX_Valid, RX_Primitive, TC1_Timeout, TC2_Timeout)
	begin
		NextState									<= State;

		TX_Primitive							<= SATA_PRIMITIVE_DIAL_TONE;

		-- general timeout
		TC1_en										<= '0';
		TC1_Load									<= '0';
		TC1_Slot									<= 0;

		-- OOB state specific timeouts
		TC2_en										<= '0';
		TC2_Load									<= '0';
		TC2_Slot									<= 0;

		HostDetected_i						<= '0';
		LinkOK_i									<= '0';
		LinkDead_i								<= '0';
		Timeout_i									<= '0';

		OOB_TX_Command_i					<= SATA_OOB_NONE;
		OOB_HandshakeComplete_i		<= '0';

		-- handle timeout with highest priority
		if (TC1_Timeout = '1') then
			TC1_en											<= '0';
			TC1_Load										<= '1';
			TC1_Slot										<= ite((SATAGeneration = SATA_GENERATION_1), TTID1_OOB_TIMEOUT_GEN1,
																		 ite((SATAGeneration = SATA_GENERATION_2), TTID1_OOB_TIMEOUT_GEN2,
																		 ite((SATAGeneration = SATA_GENERATION_3), TTID1_OOB_TIMEOUT_GEN3,
																																							 TTID1_OOB_TIMEOUT_GEN3)));
			NextState										<= ST_DEV_TIMEOUT;

		else
			case State is
				when ST_DEV_RESET =>
					-- Start automatically when Reset is deasserted.
						TC1_Load							<= '1';
						TC1_Slot							<= ite((SATAGeneration = SATA_GENERATION_1), TTID1_OOB_TIMEOUT_GEN1,
																		 ite((SATAGeneration = SATA_GENERATION_2), TTID1_OOB_TIMEOUT_GEN2,
																		 ite((SATAGeneration = SATA_GENERATION_3), TTID1_OOB_TIMEOUT_GEN3,
																																								TTID1_OOB_TIMEOUT_GEN3)));
						NextState							<= ST_DEV_WAIT_HOST_COMRESET;


				when ST_DEV_WAIT_HOST_COMRESET =>
					if (OOB_RX_Received = SATA_OOB_COMRESET) then																										-- host comreset detected
						TC1_Load							<= '1';
						TC2_Load							<= '1';
						TC1_Slot							<= ite((SATAGeneration = SATA_GENERATION_1), TTID1_OOB_TIMEOUT_GEN1,
																		 ite((SATAGeneration = SATA_GENERATION_2), TTID1_OOB_TIMEOUT_GEN2,
																		 ite((SATAGeneration = SATA_GENERATION_3), TTID1_OOB_TIMEOUT_GEN3,
																																								TTID1_OOB_TIMEOUT_GEN3)));
						TC2_Slot							<= ite((SATAGeneration = SATA_GENERATION_1), TTID2_COMRESET_TIMEOUT_GEN1,
																		 ite((SATAGeneration = SATA_GENERATION_2), TTID2_COMRESET_TIMEOUT_GEN2,
																		 ite((SATAGeneration = SATA_GENERATION_3), TTID2_COMRESET_TIMEOUT_GEN3,
																																								TTID2_COMRESET_TIMEOUT_GEN3)));
						NextState							<= ST_DEV_WAIT_AFTER_HOST_COMRESET;
						HostDetected_i 				<= '1';
					end if;

				when ST_DEV_WAIT_AFTER_HOST_COMRESET =>
					TX_Primitive						<= SATA_PRIMITIVE_DIAL_TONE;	--SATA_PRIMITIVE_ALIGN;
					TC1_en									<= '1';
					TC2_en									<= '1';

					if (OOB_RX_Received = SATA_OOB_COMRESET) then																										-- host additional comreset detected
						TC2_Load							<= '1';
						TC2_Slot							<= ite((SATAGeneration = SATA_GENERATION_1), TTID2_COMRESET_TIMEOUT_GEN1,
																		 ite((SATAGeneration = SATA_GENERATION_2), TTID2_COMRESET_TIMEOUT_GEN2,
																		 ite((SATAGeneration = SATA_GENERATION_3), TTID2_COMRESET_TIMEOUT_GEN3,
																																								TTID2_COMRESET_TIMEOUT_GEN3)));
					elsif (TC2_Timeout = '1') then
						OOB_TX_Command_i			<= SATA_OOB_COMRESET;

						NextState							<= ST_DEV_SEND_COMINIT;
					end if;

				when ST_DEV_SEND_COMINIT =>
					TX_Primitive						<= SATA_PRIMITIVE_DIAL_TONE;	--SATA_PRIMITIVE_ALIGN;
					TC1_en									<= '1';

					if (OOB_TX_Complete = '1') then
						NextState					<= ST_DEV_WAIT_HOST_COMWAKE;
					elsif ((ALLOW_STANDARD_VIOLATION = TRUE) and (OOB_RX_Received = SATA_OOB_COMWAKE)) then					-- allow premature OOB response
						NextState					<= ST_DEV_WAIT_AFTER_COMWAKE;
					end if;

				when ST_DEV_WAIT_HOST_COMWAKE =>
					TX_Primitive				<= SATA_PRIMITIVE_ALIGN;
					TC1_en							<= '1';

					if (OOB_RX_Received = SATA_OOB_COMWAKE) then																											-- host comwake detected
						TC2_Load					<= '1';
						TC2_Slot					<= ite((SATAGeneration = SATA_GENERATION_1), TTID2_COMWAKE_TIMEOUT_GEN1,
																 ite((SATAGeneration = SATA_GENERATION_2), TTID2_COMWAKE_TIMEOUT_GEN2,
																 ite((SATAGeneration = SATA_GENERATION_3), TTID2_COMWAKE_TIMEOUT_GEN3,
																																						TTID2_COMWAKE_TIMEOUT_GEN3)));
						NextState					<= ST_DEV_WAIT_AFTER_COMWAKE;
					end if;

				when ST_DEV_WAIT_AFTER_COMWAKE =>
					TC1_en							<= '1';
					TC2_en							<= '1';

					if (OOB_RX_Received = SATA_OOB_COMWAKE) then																											-- additional host cominit detected
						TC2_Load					<= '1';
						TC2_Slot					<= ite((SATAGeneration = SATA_GENERATION_1), TTID2_COMWAKE_TIMEOUT_GEN1,
																 ite((SATAGeneration = SATA_GENERATION_2), TTID2_COMWAKE_TIMEOUT_GEN2,
																 ite((SATAGeneration = SATA_GENERATION_3), TTID2_COMWAKE_TIMEOUT_GEN3,
																																						TTID2_COMWAKE_TIMEOUT_GEN3)));
					elsif (TC2_Timeout = '1') then
						OOB_TX_Command_i			<= SATA_OOB_COMWAKE;

						NextState							<= ST_DEV_SEND_COMWAKE;
					end if;

				when ST_DEV_SEND_COMWAKE =>
					TX_Primitive						<= SATA_PRIMITIVE_DIAL_TONE;	--SATA_PRIMITIVE_ALIGN;
					TC1_en									<= '1';

					if (OOB_TX_Complete = '1') then
						NextState							<= ST_DEV_OOB_HANDSHAKE_COMPLETE;
					end if;

				when ST_DEV_OOB_HANDSHAKE_COMPLETE =>
					OOB_HandshakeComplete_i	<= '1';
					TX_Primitive						<= SATA_PRIMITIVE_ALIGN;
					TC1_en 									<= '1';
					NextState								<= ST_DEV_SEND_ALIGN;

				when ST_DEV_SEND_ALIGN =>
					TX_Primitive						<= SATA_PRIMITIVE_ALIGN;
					TC1_en 									<= '1';

					if ((RX_Primitive = SATA_PRIMITIVE_ALIGN) and (RX_Valid = '1')) then												-- ALIGN detected
						NextState							<= ST_DEV_LINK_OK;
					end if;

				when ST_DEV_LINK_OK =>
					LinkOK_i								<= '1';
					TX_Primitive						<= SATA_PRIMITIVE_NONE;

					if (OOB_RX_Received /= SATA_OOB_NONE) then
						NextState							<= ST_DEV_LINK_DEAD;
					end if;

				when ST_DEV_LINK_DEAD =>
					-- Reset must be asserted to leave this state.
					LinkDead_i							<= '1';

						TC1_Load							<= '1';
						TC1_Slot							<= ite((SATAGeneration = SATA_GENERATION_1), TTID1_OOB_TIMEOUT_GEN1,
																		 ite((SATAGeneration = SATA_GENERATION_2), TTID1_OOB_TIMEOUT_GEN2,
																		 ite((SATAGeneration = SATA_GENERATION_3), TTID1_OOB_TIMEOUT_GEN3,
																																							 TTID1_OOB_TIMEOUT_GEN3)));
						NextState							<= ST_DEV_WAIT_HOST_COMRESET;

				when ST_DEV_TIMEOUT =>
					-- Reset must be asserted to leave this state.
					Timeout_i								<= '1';

						TC1_Load							<= '1';
						TC1_Slot							<= ite((SATAGeneration = SATA_GENERATION_1), TTID1_OOB_TIMEOUT_GEN1,
																		 ite((SATAGeneration = SATA_GENERATION_2), TTID1_OOB_TIMEOUT_GEN2,
																		 ite((SATAGeneration = SATA_GENERATION_3), TTID1_OOB_TIMEOUT_GEN3,
																																							 TTID1_OOB_TIMEOUT_GEN3)));
						NextState							<= ST_DEV_WAIT_HOST_COMRESET;

			end case;
		end if;
	end process;

	HostDetected						<= HostDetected_i;
	LinkOK									<= LinkOK_i;
	LinkDead								<= LinkDead_i;
	Timeout									<= Timeout_i;

	OOB_TX_Command					<= OOB_TX_Command_i;
	OOB_HandshakeComplete		<= OOB_HandshakeComplete_i;


	-- overall timeout counter
	TC1 : entity PoC.io_TimingCounter
		generic map (							-- timing table
			TIMING_TABLE				=> TC1_TIMING_TABLE
		)
		port map (
			Clock								=> Clock,
			Enable							=> TC1_en,
			Load								=> TC1_Load,
			Slot								=> TC1_Slot,
			Timeout							=> TC1_Timeout
		);

	-- timeout counter for *_WAIT_AFTER_* states
	TC2 : entity PoC.io_TimingCounter
		generic map (							-- timing table
			TIMING_TABLE				=> TC2_TIMING_TABLE
		)
		port map (
			Clock								=> Clock,
			Enable							=> TC2_en,
			Load								=> TC2_Load,
			Slot								=> TC2_Slot,
			Timeout							=> TC2_Timeout
		);

	-- debug port
	-- ===========================================================================
	genDebugPort : if (ENABLE_DEBUGPORT = TRUE) generate
		function dbg_EncodeState(st : T_STATE) return std_logic_vector is
		begin
			return to_slv(T_STATE'pos(st), log2ceilnz(T_STATE'pos(T_STATE'high) + 1));
		end function;

		function dbg_GenerateEncodings return string is
			variable  l : STD.TextIO.line;
		begin
			for i in T_STATE loop
				STD.TextIO.write(l, str_replace(T_STATE'image(i), "st_dev_", ""));
				STD.TextIO.write(l, ';');
			end loop;
			return  l.all;
		end function;

--		constant dummy : boolean := dbg_ExportEncoding("OOBControl (Device)", dbg_GenerateEncodings,  PROJECT_DIR & "ChipScope/TokenFiles/FSM_OOBControl_Device.tok");
	begin
		DebugPortOut.FSM												<= dbg_EncodeState(State);
		DebugPortOut.DeviceOrHostDetected				<= HostDetected_i;
		DebugPortOut.Timeout										<= Timeout_i;
		DebugPortOut.LinkOK											<= LinkOK_i;
		DebugPortOut.LinkDead										<= LinkDead_i;

		DebugPortOut.OOB_TX_Command							<= OOB_TX_Command_i;
		DebugPortOut.OOB_TX_Complete						<= OOB_TX_Complete;
		DebugPortOut.OOB_RX_Received						<= OOB_RX_Received;
		DebugPortOut.OOB_HandshakeComplete			<= OOB_HandshakeComplete_i;
	end generate;
end;
