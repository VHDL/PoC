LIBRARY IEEE;
USE			IEEE.STD_LOGIC_1164.ALL;
USE			IEEE.NUMERIC_STD.ALL;

LIBRARY PoC;
USE			PoC.utils.ALL;
USE			PoC.vectors.ALL;
USE			PoC.lcd.ALL;


ENTITY lcd_LCDSynchronizer IS
	GENERIC (
		CLOCK_FREQ_MHZ			: REAL		:= 100.0			-- 100 MHz
	);
	PORT (
		Clock								: IN	STD_LOGIC;
		Reset								: IN	STD_LOGIC;
		
		Synchronize					: IN	STD_LOGIC;
		Synchronized				: OUT	STD_LOGIC;
		
		Column							: OUT	T_LCD_COLUMN_INDEX;
		Row									:	OUT	T_LCD_ROW_INDEX;
		Char								: IN	T_LCD_CHAR;
		
		-- LCD interface
		LCD_en							:	OUT	STD_LOGIC;
		LCD_rw							: OUT	STD_LOGIC;
		LCD_rs							: OUT	STD_LOGIC;								-- LCD Register Select
		LCD_Data_o					: OUT	T_SLV_4;
    LCD_Data_t    			: OUT STD_LOGIC;
    LCD_Data_i    			: IN  T_SLV_4
	);
END;


ARCHITECTURE rtl OF lcd_LCDSynchronizer IS
	ATTRIBUTE KEEP		: STRING;

	TYPE T_STATE IS (
		ST_RESET,
		ST_INIT_SET_FUNCTION, ST_INIT_SET_FUNCTION_WAIT,
		ST_INIT_DISPLAY_ON, ST_INIT_DISPLAY_ON_WAIT,
		ST_INIT_DISPLAY_CLEAR, ST_INIT_DISPLAY_CLEAR_WAIT,
		ST_INIT_ENTRY_MODE, ST_INIT_ENTRY_MODE_WAIT,
		ST_IDLE,
		ST_GO_HOME, ST_GO_HOME_WAIT,
		ST_WRITE_CHAR, ST_WRITE_CHAR_WAIT,
		ST_FINISHED
	);
		
	SIGNAL State			: T_STATE			:= ST_RESET;
	SIGNAL NextState	: T_STATE;

	CONSTANT COLAC_BW				: POSITIVE																			:= T_LCD_COLUMN_INDEX_BW;
	CONSTANT ROWAC_BW				: POSITIVE																			:= T_LCD_ROW_INDEX_BW;

	SIGNAL ColAC_inc				: STD_LOGIC;
	SIGNAL ColAC_Load				: STD_LOGIC;
	SIGNAL ColAC_Address		: STD_LOGIC_VECTOR(COLAC_BW - 1 DOWNTO 0);
	SIGNAL ColAC_Address_us	: UNSIGNED(COLAC_BW - 1 DOWNTO 0);
	SIGNAL ColAC_Finished		: STD_LOGIC;

	SIGNAL RowAC_inc				: STD_LOGIC;
	SIGNAL RowAC_Load				: STD_LOGIC;
	SIGNAL RowAC_Address		: STD_LOGIC_VECTOR(ROWAC_BW - 1 DOWNTO 0);
	SIGNAL RowAC_Address_us	: UNSIGNED(ROWAC_BW - 1 DOWNTO 0);
	SIGNAL RowAC_Finished		: STD_LOGIC;

	SIGNAL LCDI_Strobe			: STD_LOGIC;
	SIGNAL LCDI_Address			: STD_LOGIC;
	SIGNAL LCDI_Data				: T_SLV_8;
	SIGNAL LCDI_Ready				: STD_LOGIC;

	SIGNAL CSP_Trigger_1		: STD_LOGIC;
	ATTRIBUTE KEEP OF CSP_Trigger_1 : SIGNAL IS "TRUE";

BEGIN

	PROCESS(Clock)
	BEGIN
		IF rising_edge(Clock) THEN
			IF (Reset = '1') THEN
				State		<= ST_RESET;
			ELSE
				State		<= NextState;
			END IF;
		END IF;
	END PROCESS;
	
	
	PROCESS(State, LCDI_Ready, Synchronize, Char, RowAC_Address_us, ColAC_Finished, RowAC_Finished)
	BEGIN
		NextState					<= State;
		
		Synchronized			<= '0';
		
		ColAC_inc					<= '0';
		ColAC_Load				<= '0';
		RowAC_inc					<= '0';
		RowAC_Load				<= '0';
		
		LCDI_Strobe				<= '0';
		LCDI_Address			<= '0';
		LCDI_Data					<= LCDCMD_NONE;
		
		CSP_Trigger_1			<= '0';
		
		CASE State IS
			WHEN ST_RESET =>
				IF (LCDI_Ready = '1') THEN
					CSP_Trigger_1	<= '1';
					
					NextState			<= ST_INIT_SET_FUNCTION;
				END IF;
	
			WHEN ST_INIT_SET_FUNCTION =>
				LCDI_Strobe			<= '1';
				LCDI_Address		<= '0';
				LCDI_Data				<= LCDCMD_SET_FUNCTION;
				
				NextState				<= ST_INIT_SET_FUNCTION_WAIT;
			
			WHEN ST_INIT_SET_FUNCTION_WAIT =>
				IF (LCDI_Ready = '1') THEN
					NextState			<= ST_INIT_DISPLAY_ON;
				END IF;
			
			WHEN ST_INIT_DISPLAY_ON =>
				LCDI_Strobe			<= '1';
				LCDI_Address		<= '0';
				LCDI_Data				<= lcd_display_on(FALSE, FALSE);
				
				NextState				<= ST_INIT_DISPLAY_ON_WAIT;
			
			WHEN ST_INIT_DISPLAY_ON_WAIT =>
				IF (LCDI_Ready = '1') THEN
					NextState			<= ST_INIT_DISPLAY_CLEAR;
				END IF;
			
			WHEN ST_INIT_DISPLAY_CLEAR =>
				LCDI_Strobe			<= '1';
				LCDI_Address		<= '0';
				LCDI_Data				<= LCDCMD_DISPLAY_CLEAR;
				
				NextState				<= ST_INIT_DISPLAY_CLEAR_WAIT;
			
			WHEN ST_INIT_DISPLAY_CLEAR_WAIT =>
				IF (LCDI_Ready = '1') THEN
					NextState			<= ST_INIT_ENTRY_MODE;
				END IF;
			
			WHEN ST_INIT_ENTRY_MODE =>
				LCDI_Strobe			<= '1';
				LCDI_Address		<= '0';
				LCDI_Data				<= LCDCMD_ENTRY_MODE;
				
				NextState				<= ST_INIT_ENTRY_MODE_WAIT;
			
			WHEN ST_INIT_ENTRY_MODE_WAIT =>
				IF (LCDI_Ready = '1') THEN
					NextState			<= ST_IDLE;
				END IF;
			
			WHEN ST_IDLE =>
				IF (Synchronize = '1') THEN
					ColAC_Load			<= '1';
					RowAC_Load			<= '1';

					NextState			<= ST_GO_HOME;
				END IF;
			
			WHEN ST_GO_HOME =>
				LCDI_Strobe			<= '1';
				LCDI_Address		<= '0';
				LCDI_Data				<= lcd_go_home(RowAC_Address_us);
				
				NextState				<= ST_GO_HOME_WAIT;
			
			WHEN ST_GO_HOME_WAIT =>
				IF (LCDI_Ready = '1') THEN
					NextState			<= ST_WRITE_CHAR;
				END IF;
	
			WHEN ST_WRITE_CHAR =>
				ColAC_inc				<= '1';
			
				LCDI_Strobe			<= '1';
				LCDI_Address		<= '1';
				LCDI_Data				<= LCD_Char2Bin(Char);
				
				NextState				<= ST_WRITE_CHAR_WAIT;
			
			WHEN ST_WRITE_CHAR_WAIT =>
				IF (LCDI_Ready = '1') THEN
					IF (ColAC_Finished = '1') THEN
						IF (RowAC_Finished = '1') THEN
							ColAC_Load	<= '1';
							RowAC_Load	<= '1';
							
							NextState		<= ST_FINISHED;
						ELSE
							ColAC_Load	<= '1';
							RowAC_inc		<= '1';
				
							NextState		<= ST_GO_HOME;
						END IF;
					ELSE
						NextState			<= ST_WRITE_CHAR;
					END IF;
				END IF;
	
			WHEN ST_FINISHED =>
				Synchronized			<= '1';
				
				NextState					<= ST_IDLE;
	
		END CASE;
	END PROCESS;

	ColAC : ENTITY L_Global.AddressCounter
		GENERIC MAP (
			COUNTER_BW					=> COLAC_BW
		)
		PORT MAP (
			Clock								=> Clock,																							-- clock
			inc									=> ColAC_inc,																					-- enable counter
			Load								=> ColAC_Load,																				-- load start and forward input
			Address_Start				=> to_slv(0, COLAC_BW),																-- start address
			Address_Step				=> to_slv(1, COLAC_BW),																-- step between two addresses
			Address_End					=> to_slv(MAX_LCD_COLUMN_COUNT, COLAC_BW),						-- end address

			Address							=> ColAC_Address,																			-- currend address
			Counter_Finished		=> ColAC_Finished																			-- active if end address is reached
		);

	RowAC : ENTITY L_Global.AddressCounter
		GENERIC MAP (
			COUNTER_BW					=> ROWAC_BW
		)
		PORT MAP (
			Clock								=> Clock,																							-- clock
			inc									=> RowAC_inc,																					-- enable counter
			Load								=> RowAC_Load,																				-- load start and forward input
			Address_Start				=> to_slv(0, ROWAC_BW),																-- start address
			Address_Step				=> to_slv(1, ROWAC_BW),																-- step between two addresses
			Address_End					=> to_slv(MAX_LCD_ROW_COUNT - 1, ROWAC_BW),						-- end address

			Address							=> RowAC_Address,																			-- currend address
			Counter_Finished		=> RowAC_Finished																			-- active if end address is reached
		);

	ColAC_Address_us	<= unsigned(ColAC_Address);
	RowAC_Address_us	<= unsigned(RowAC_Address);

	Column	<= to_integer(ColAC_Address_us);
	Row			<= to_integer(RowAC_Address_us);

	LCDInterface : ENTITY L_LCD.lcd4
		PORT MAP (
			-- Global Reset and Clock
			clk					=> Clock,
			rst					=> Reset,

			-- Upper Layer Interface
			stb      		=> LCDI_Strobe,
			addr     		=> LCDI_Address,
			din      		=> LCDI_Data,
			rdy      		=> LCDI_Ready,
			
			-- LCD Connections
			lcd_e   		=> LCD_en,
			lcd_rs  		=> LCD_rs,
			lcd_rw  		=> LCD_rw,
			lcd_dat_o 	=> LCD_Data_o,
			lcd_dat_t 	=> LCD_Data_t,
			lcd_dat_i	  => LCD_Data_i
		);
END;
