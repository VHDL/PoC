-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- 
-- ============================================================================
-- Authors:					Martin Zabel
--									Patrick Lehmann
-- 
-- Module:					Instantiates Chip-Specific DDR Output Registers for Xilinx FPGAs.
--
-- Description:
-- ------------------------------------
--		See PoC.io.ddrio.out for interface description.
--		
-- License:
-- ============================================================================
-- Copyright 2007-2015 Technische Universitaet Dresden - Germany,
--										 Chair for VLSI-Design, Diagnostics and Architecture
-- 
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
-- 
--		http://www.apache.org/licenses/LICENSE-2.0
-- 
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- ============================================================================


library IEEE;
use			IEEE.std_logic_1164.ALL;

library	UniSim;
use			UniSim.vComponents.all;


entity ddrio_out_xilinx is
	generic (
		NO_OE				: boolean		:= false;
		INIT_VALUE	: BIT				:= '1';
		WIDTH				: positive
	);
	port (
		clk		: in	std_logic;
		ce		: in	std_logic;
		dh		: in	std_logic_vector(WIDTH-1 downto 0);
		dl		: in	std_logic_vector(WIDTH-1 downto 0);
		oe		: in	std_logic;
		q			: out	std_logic_vector(WIDTH-1 downto 0)
	);
end entity;


architecture rtl of ddrio_out_xilinx is

begin
	gen : for i in 0 to WIDTH - 1 generate
		signal o : std_logic;
	begin
		dff : ODDR
			generic map(
				DDR_CLK_EDGE	=> "SAME_EDGE",
				INIT					=> INIT,
				SRTYPE				=> "SYNC"
			)
			port map (
				Q		=> o,
				C		=> clk,
				CE	=> ce,
				D1	=> dh(i),
				D2	=> dl(i),
				R		=> '0',
				S		=> '0'
			);

		genOE : if not NO_OE generate
			signal oe_n : std_logic;
			signal t    : std_logic;
		 begin
			oe_n <= not oe;
			 
			oeff : ODDR
				generic map(
					DDR_CLK_EDGE	=> "SAME_EDGE",
					INIT					=> '1',
					SRTYPE				=> "SYNC"
				)
				port map (
					Q		=> t,
					C		=> clk,
					CE	=> ce,
					D1	=> oe_n,
					D2	=> oe_n,
					R		=> '0',
					S		=> '0'
				);

			q(i) <= o when t = '0' else 'Z';  -- 't' is low-active!
		end generate genOE;

		genNoOE : if NO_OE generate
			q(i) <= o;
		end generate genNoOE;
	end generate;
end architecture;
