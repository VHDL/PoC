-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- =============================================================================
-- Authors:					G. Martin
--
-- Entity:					arith_counter_bcd_TestHarness
--
-- Description:
-- -------------------------------------
-- Test harness for arith_counter_bcd
--
-- License:
-- =============================================================================
-- Copyright 2025-2025 The PoC-Library Authors
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--		http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- =============================================================================

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library osvvm;
context osvvm.OsvvmContext;

library PoC;
use PoC.utils.all;
use PoC.strings.all;
use PoC.physical.all;

entity arith_counter_bcd_TestHarness is
end entity;

architecture TestHarness of arith_counter_bcd_TestHarness is
  constant TPERIOD_CLOCK : time := 10 ns;
  constant CLOCK_FREQ : FREQ := 100 MHz;
  constant DIGITS : positive := 3;

  signal Clock : std_logic := '1';
  signal Reset : std_logic := '1';
  signal Reset_aux : std_logic := '0';
  signal inc : std_logic := '0';
  signal Value : T_BCD_VECTOR(DIGITS - 1 downto 0);

  component arith_counter_bcd_TestController is
    generic (
      DIGITS : positive := 3
    );
    port (
      Clock     : in std_logic;
      Reset     : in std_logic;
      Reset_aux : out std_logic;
      inc       : out std_logic;
      Value     : in T_BCD_VECTOR(DIGITS - 1 downto 0)
    );
  end component;

begin

  Osvvm.ClockResetPkg.CreateClock(
    Clk    => Clock, 
    Period => TPERIOD_CLOCK
  );

  Osvvm.ClockResetPkg.CreateReset(
    Reset       => Reset, 
    ResetActive => '1', 
    Clk         => Clock, 
    Period      => 5 * TPERIOD_CLOCK, 
    tpd         => 0 ns
  );

  UUT: entity PoC.arith_counter_bcd
    generic map (
      DIGITS => DIGITS
    )
    port map (
      clk => Clock,
      rst => Reset or Reset_aux,
      inc => inc,
      val => Value
    );
    
  TestCtrl: component arith_counter_bcd_TestController
    generic map (
      DIGITS => DIGITS
    )
    port map (
      Clock     => Clock,
      Reset     => Reset,
      Reset_aux => Reset_aux,
      inc       => inc,
      Value     => Value
    );
end architecture;