

package misc is

end package;

package body misc is

end package body;
