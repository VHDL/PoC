-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
--
-- =============================================================================
-- Authors:					Patrick Lehmann
--
-- Module:					Primtive Detector for SATA Link Layer
--
-- Description:
-- ------------------------------------
-- Detects primitives in the incoming data stream from the physical link. If
-- a primitive X is continued via the CONT primitive and scrambled dummy data,
-- this unit outputs X continously until a new primitve (except ALIGN) arrives.
--
-- License:
-- =============================================================================
-- Copyright 2007-2015 Technische Universitaet Dresden - Germany
--										 Chair for VLSI-Design, Diagnostics and Architecture
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--		http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- =============================================================================

LIBRARY IEEE;
USE			IEEE.STD_LOGIC_1164.ALL;
USE			IEEE.NUMERIC_STD.ALL;

LIBRARY PoC;
USE			PoC.utils.ALL;
USE			PoC.vectors.ALL;
USE			PoC.components.ALL;
USE			PoC.sata.ALL;


ENTITY sata_PrimitiveDetector IS
	PORT (
		Clock									: IN	STD_LOGIC;

		RX_DataIn							: IN	T_SLV_32;
		RX_CharIsK						: IN	T_SLV_4;

		Primitive							: OUT	T_SATA_PRIMITIVE
	);
END;

-- Example waveform
-- """"""""""""""""""""""
-- Primitive_i							< TX_RDY ><  CONT  ><  XXXX  ><  XXXX  >< RX_RDY ><  CONT  ><  XXXX  ><  XXXX  >
-- PrimitiveReg_ctrl_rst		__________""""""""""______________________________""""""""""____________________
-- PrimitiveReg_ctrl_set		""""""""""______________________________""""""""""______________________________
-- PrimitiveReg_ctrl				""""""""""""""""""""______________________________""""""""""____________________
-- PrimitiveReg_en					""""""""""______________________________""""""""""______________________________
-- PrimitiveReg_d						<  ????  >< TX_RDY >< TX_RDY >< TX_RDY >< TX_RDY >< RX_RDY >< RX_RDY >< RX_RDY >
-- Primitive								< TX_RDY >< TX_RDY >< TX_RDY >< TX_RDY >< RX_RDY >< RX_RDY >< RX_RDY >< RX_RDY >

ARCHITECTURE rtl OF sata_PrimitiveDetector IS
	SIGNAL Primitive_i							: T_SATA_PRIMITIVE;

	SIGNAL PrimitiveReg_ctrl_rst		: STD_LOGIC;
	SIGNAL PrimitiveReg_ctrl_set		: STD_LOGIC;
	SIGNAL PrimitiveReg_ctrl				: STD_LOGIC						:= '1';
	SIGNAL PrimitiveReg_en					: STD_LOGIC;
	SIGNAL PrimitiveReg_d						: T_SATA_PRIMITIVE		:= SATA_PRIMITIVE_NONE;

BEGIN
	Primitive_i		<= to_sata_primitive(RX_DataIn, RX_CharIsK);

	-- ===========================================================================
	-- SATA_PRIMITIVE_CONT feature
	-- ===========================================================================
	-- PrimitiveReg_ctrl - if CONT ocours -> disable PrimitiveReg
	PrimitiveReg_ctrl_rst		<= to_sl(Primitive_i = SATA_PRIMITIVE_CONT);
	PrimitiveReg_ctrl_set		<= NOT to_sl((Primitive_i = SATA_PRIMITIVE_CONT) OR
																			 (Primitive_i = SATA_PRIMITIVE_ALIGN) OR
																			 (Primitive_i = SATA_PRIMITIVE_NONE) OR
																			 (Primitive_i = SATA_PRIMITIVE_ILLEGAL));

	PrimitiveReg_ctrl	<= ffsr(q => PrimitiveReg_ctrl, rst => PrimitiveReg_ctrl_rst, set => PrimitiveReg_ctrl_set) WHEN rising_edge(Clock);
	PrimitiveReg_en		<= (PrimitiveReg_ctrl OR PrimitiveReg_ctrl_set) AND NOT PrimitiveReg_ctrl_rst;

	-- PrimitiveReg - save last received primitive
	PROCESS(Clock)
	BEGIN
		IF rising_edge(Clock) THEN
			IF (PrimitiveReg_en = '1') AND NOT (Primitive_i = SATA_PRIMITIVE_ALIGN) THEN
				PrimitiveReg_d	<= Primitive_i;
			END IF;
		END IF;
	END PROCESS;

	Primitive	<= Primitive_i WHEN (PrimitiveReg_en = '1') ELSE PrimitiveReg_d;
END;
