LIBRARY IEEE;
USE			IEEE.STD_LOGIC_1164.ALL;
USE			IEEE.NUMERIC_STD.ALL;

LIBRARY PoC;
USE			PoC.functions.ALL;

-- Usage
-- ====================================
 --LIBRARY	L_SATAController;
 --USE			L_SATAController.SATATransceiverTypes.ALL;

PACKAGE SATATransceiverTypes IS
	TYPE T_SATA_TRANSCEIVER_COMMON_SIGNALS IS RECORD
		RefClockIn_75_MHz			: STD_LOGIC;
		RefClockIn_150_MHz		: STD_LOGIC;
	END RECORD;

	TYPE T_SATA_TRANSCEIVER_PRIVATE_SIGNALS IS RECORD
		TX_n									: STD_LOGIC;
		TX_p									: STD_LOGIC;
		RX_n									: STD_LOGIC;
		RX_p									: STD_LOGIC;
	END RECORD;
	
	TYPE T_SATA_TRANSCEIVER_PRIVATE_SIGNALS_VECTOR IS ARRAY(NATURAL RANGE <>) OF T_SATA_TRANSCEIVER_PRIVATE_SIGNALS;
END SATATransceiverTypes;

PACKAGE BODY SATATransceiverTypes IS

END PACKAGE BODY;
