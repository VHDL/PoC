-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- ============================================================================
-- Authors:					Patrick Lehmann
--
-- Context:					Provides all packages from <PoCRoot>/src/common.
--
-- Description:
-- ------------------------------------
--		This package provides all common packages as a single context.
--
-- License:
-- ============================================================================
-- Copyright 2007-2015 Technische Universitaet Dresden - Germany,
--										 Chair for VLSI-Design, Diagnostics and Architecture
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--		http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- ============================================================================

context Common is
	library PoC ;
	use PoC.config.all;
	use PoC.debug.all;
	use PoC.FileIO.all;
	use PoC.math.all;
	use PoC.physical.all;
	use PoC.strings.all;
	use PoC.utils.all;
	use PoC.vectors.all;
end context;
