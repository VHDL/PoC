-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- =============================================================================
-- Authors:					Gustavo Martin
--
-- Entity:					arith_trng_TestController
--
-- Description:
-- -------------------------------------
-- Simple test for arith_trng component (True Random Number Generator)
--
-- License:
-- =============================================================================
-- Copyright 2025-2025 The PoC-Library Authors
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--		http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- =============================================================================

library IEEE;
use     IEEE.std_logic_1164.all;
use     IEEE.numeric_std.all;

library osvvm;
context osvvm.OsvvmContext;

library PoC;
use     PoC.utils.all;

architecture Simple of arith_trng_TestController is
	signal TestDone : integer_barrier := 1;

	constant TCID : AlertLogIDType :=  NewID("TestCtrl");

begin
	ControlProc: process
		constant ProcID : AlertLogIDType := NewID("ControlProc", TCID);
		constant TIMEOUT : time := 10 ms;
	begin
		SetTestName("arith_trng_Simple");

		SetLogEnable(PASSED, FALSE);
		SetLogEnable(INFO,   FALSE);
		SetLogEnable(DEBUG,  FALSE);
		wait for 0 ns; wait for 0 ns;

		TranscriptOpen;
		SetTranscriptMirror(TRUE);

		wait until Reset = '0';
		ClearAlerts;

		WaitForBarrier(TestDone, TIMEOUT);
		AlertIf(ProcID, now >= TIMEOUT,     "Test finished due to timeout");
		AlertIf(ProcID, GetAffirmCount < 1, "Test is not Self-Checking");

		EndOfTestReports(ReportAll => TRUE);
		std.env.stop;
	end process;

	CheckerProc: process
		constant ProcID : AlertLogIDType := NewID("CheckerProc", TCID);
		constant NUM_SAMPLES : natural := 100;
		
		variable prev_rnd : std_logic_vector(rnd'range);
		variable changes : natural := 0;
		variable has_zeros : boolean := false;
		variable has_ones : boolean := false;
	begin
		wait until Reset = '0';
		WaitForClock(Clock);

		-- NOTE: TRNGs rely on hardware phenomena (metastability, jitter, etc.) that
		-- are not accurately modeled in simulation. This test verifies basic functionality
		-- but cannot validate true randomness. True TRNG validation must be done on
		-- actual hardware using tools like dieharder.
		
		-- Verify the component produces output
		prev_rnd := rnd;
		WaitForClock(Clock);
		
		-- Sample multiple times to check if any variation occurs
		for i in 1 to NUM_SAMPLES loop
			if rnd /= prev_rnd then
				changes := changes + 1;
			end if;
			-- Check for bit patterns
			if rnd = (rnd'range => '0') then
				has_zeros := true;
			end if;
			if rnd = (rnd'range => '1') then
				has_ones := true;
			end if;
			prev_rnd := rnd;
			WaitForClock(Clock);
		end loop;

		-- Basic sanity checks that are simulation-friendly
		-- Note: In simulation, TRNG may produce constant or deterministic output
		Log(ProcID, "TRNG changes observed: " & integer'image(changes) & 
			" out of " & integer'image(NUM_SAMPLES) & " samples", INFO);
		
		-- Check that the output is defined (not 'U' or 'X')
		AffirmIf(ProcID, not is_x(rnd), "TRNG output should be defined (not X or U)");

		-- Verify component can be read without errors
		for i in 1 to 10 loop
			WaitForClock(Clock);
			AffirmIf(ProcID, not is_x(rnd), "TRNG continues to produce defined output");
		end loop;

		-- Note to user: Actual randomness verification must be done on hardware
		Log(ProcID, "WARNING: TRNG randomness cannot be verified in simulation.", WARNING);
		Log(ProcID, "Verify randomness on target hardware using dieharder or similar tools.", WARNING);

		WaitForBarrier(TestDone);
		wait;
	end process;
end architecture;

configuration arith_trng_Simple of arith_trng_TestHarness is
	for TestHarness
		for TestCtrl: arith_trng_TestController
			use entity work.arith_trng_TestController(Simple);
		end for;
	end for;
end configuration;
