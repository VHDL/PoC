-- EMACS settings: -*-  tab-width:2  -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- 
-- ============================================================================================================================================================
-- Description:     Project specific configuration.
--                  This is a template file. 
--                  The global package common/config evaluates the settings declared in this file.
--
-- Usage:
--                  1) Copy this file into your project's source directory and rename it to my_config.vhdl.
--                  2) Add file to library "poc" in your synthesis tool.
--                  3) Change setup appropriately.
--
-- Authors:         Thomas B. Preusser
--                  Martin Zabel
--                  Patrick Lehmann
-- ============================================================================================================================================================
-- Copyright 2007-2013 Technische Universität Dresden - Germany, Chair for VLSI-Design, Diagnostics and Architecture
-- 
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
-- 
--    http://www.apache.org/licenses/LICENSE-2.0
-- 
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- ============================================================================================================================================================
library PoC;

package my_config is
  -- Change these lines to setup configuration.
  constant MY_DEVICE : string := "XC5VLX50T"; -- e.g. XC5VLX50T, EP2SGX90
 
end my_config;

package body my_config is

end my_config;

