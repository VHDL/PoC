LIBRARY IEEE;
USE			IEEE.STD_LOGIC_1164.ALL;
USE			IEEE.NUMERIC_STD.ALL;

LIBRARY PoC;
USE			PoC.functions.ALL;

-- Usage
-- ====================================
 --LIBRARY	L_SATAController;
 --USE			L_SATAController.SATATransceiverTypes.ALL;

PACKAGE SATATransceiverTypes IS
	TYPE T_SATA_TRANSCEIVER_COMMON_IN_SIGNALS IS RECORD
		RefClockIn_150_MHz		: STD_LOGIC;
	END RECORD;

	TYPE T_SATA_TRANSCEIVER_PRIVATE_IN_SIGNALS IS RECORD
		RX_n									: STD_LOGIC;
		RX_p									: STD_LOGIC;
	END RECORD;
	TYPE T_SATA_TRANSCEIVER_PRIVATE_OUT_SIGNALS IS RECORD
		TX_n									: STD_LOGIC;
		TX_p									: STD_LOGIC;
	END RECORD;
	
	TYPE T_SATA_TRANSCEIVER_COMMON_IN_SIGNALS_VECTOR		IS ARRAY(NATURAL RANGE <>) OF T_SATA_TRANSCEIVER_COMMON_IN_SIGNALS;
	TYPE T_SATA_TRANSCEIVER_PRIVATE_IN_SIGNALS_VECTOR		IS ARRAY(NATURAL RANGE <>) OF T_SATA_TRANSCEIVER_PRIVATE_IN_SIGNALS;
	TYPE T_SATA_TRANSCEIVER_PRIVATE_OUT_SIGNALS_VECTOR	IS ARRAY(NATURAL RANGE <>) OF T_SATA_TRANSCEIVER_PRIVATE_OUT_SIGNALS;
	
END SATATransceiverTypes;

PACKAGE BODY SATATransceiverTypes IS

END PACKAGE BODY;
