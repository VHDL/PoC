-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- =============================================================================
-- Authors:					Patrick Lehmann
-- 									Martin Zabel
--
-- Entity:					FIS Decoder for SATA Transport Layer
--
-- Description:
-- -------------------------------------
-- See notes on module 'sata_TransportLayer'.
--
-- License:
-- =============================================================================
-- Copyright 2007-2015 Technische Universitaet Dresden - Germany
--										 Chair for VLSI-Design, Diagnostics and Architecture
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--		http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- =============================================================================

library IEEE;
use			IEEE.STD_LOGIC_1164.all;
use			IEEE.NUMERIC_STD.all;

library PoC;
use			PoC.config.all;
use			PoC.utils.all;
use			PoC.vectors.all;
use			PoC.strings.all;
use			PoC.debug.all;
use			PoC.sata.all;
use			PoC.satadbg.all;


entity sata_FISDecoder is
	generic (
		DEBUG													: boolean						:= FALSE;
		ENABLE_DEBUGPORT							: boolean						:= FALSE
	);
	port (
		Clock													: in	std_logic;
		Reset													: in	std_logic;

		Status												: out	T_SATA_FISDECODER_STATUS;
		FISType												: out T_SATA_FISTYPE;
		UpdateATARegisters						: out	std_logic;
		ATADeviceRegisters						: out	T_SATA_ATA_DEVICE_REGISTERS;

		-- debugPort
		DebugPortOut									: out	T_SATADBG_TRANS_FISD_OUT;

		-- TransportLayer RX_ interface
		RX_Valid											: out	std_logic;
		RX_Data												: out	T_SLV_32;
		RX_SOP												: out	std_logic;
		RX_EOP												: out	std_logic;
		RX_Ack												: in	std_logic;

		-- LinkLayer CSE
		Link_Status										: in	T_SATA_LINK_STATUS;

		-- LinkLayer FIFO interface
		Link_RX_Ack										: out	std_logic;
		Link_RX_Data									: in	T_SLV_32;
		Link_RX_SOF										: in	std_logic;
		Link_RX_EOF										: in	std_logic;
		Link_RX_Valid									: in	std_logic;

		-- LinkLayer FS-FIFO interface
		Link_RX_FS_Ack								: out	std_logic;
		Link_RX_FS_CRCOK							: in	std_logic;
		Link_RX_FS_SyncEsc						: in	std_logic;
		Link_RX_FS_Valid							: in	std_logic
	);
end entity;


architecture rtl of sata_FISDecoder is
	attribute KEEP									: boolean;
	attribute FSM_ENCODING					: string;

	type T_STATE is (
		ST_RESET, ST_IDLE, ST_CHECK_FISTYPE,
		ST_FIS_REG_DEV_HOST_WORD_1,	ST_FIS_REG_DEV_HOST_WORD_2,	ST_FIS_REG_DEV_HOST_WORD_3,	ST_FIS_REG_DEV_HOST_WORD_4,
		ST_FIS_PIO_SETUP_WORD_1,		ST_FIS_PIO_SETUP_WORD_2,		ST_FIS_PIO_SETUP_WORD_3,		ST_FIS_PIO_SETUP_WORD_4,
		ST_FIS_DATA_1,							ST_FIS_DATA_N,
		ST_RECEIVE_OK, ST_STATUS_ERROR, ST_STATUS_CRC_ERROR,
		ST_DISCARD_FRAME_1, ST_DISCARD_FRAME_N
	);

	-- alias-Definitions for FISType Register Transfer Device => Host (34h)
	-- ====================================================================================
	-- Word 0
	alias Alias_FISType										: T_SLV_8													is Link_RX_Data(7 downto 0);
	alias Alias_FlagReg										: T_SLV_8													is Link_RX_Data(15 downto 8);				-- Flag bits
	alias Alias_StatusReg									: T_SLV_8													is Link_RX_Data(23 downto 16);			-- Status register
	alias Alias_ErrorReg									: T_SLV_8													is Link_RX_Data(31 downto 24);			-- Error register
	-- Word 1
	alias Alias_LBA0											: T_SLV_8													is Link_RX_Data(7 downto 0);				-- Sector Number
	alias Alias_LBA16											: T_SLV_8													is Link_RX_Data(15 downto 8);				-- Cylinder Low
	alias Alias_LBA32											: T_SLV_8													is Link_RX_Data(23 downto 16);			-- Cylinder High
	alias Alias_Head											: T_SLV_4													is Link_RX_Data(27 downto 24);			-- Head number
	alias Alias_Device										: std_logic_vector(0 downto 0)		is Link_RX_Data(28 downto 28);			-- Device number

	-- Word 2
	alias Alias_LBA8											: T_SLV_8													is Link_RX_Data(7 downto 0);				-- Sector Number expanded
	alias Alias_LBA24											: T_SLV_8													is Link_RX_Data(15 downto 8);				-- Cylinder Low expanded
	alias Alias_LBA40											: T_SLV_8													is Link_RX_Data(23 downto 16);			-- Cylinder High expanded

	-- Word 3
	alias Alias_SecCount0									: T_SLV_8													is Link_RX_Data(7 downto 0);				-- Sector Count
	alias Alias_SecCount8									: T_SLV_8													is Link_RX_Data(15 downto 8);				-- Sector Count expanded

	-- Word 4
	alias Alias_TransferCount							: T_SLV_16												is Link_RX_Data(15 downto 0);				-- Transfer Count

	-- alias-Definitions for FISType PIO Setup (5Fh)
	-- ====================================================================================
	-- Word 3
	alias Alias_EndStatusReg							: T_SLV_8													is Link_RX_Data(31 downto 24);			-- EndStatus Register

	signal State													: T_STATE													:= ST_RESET;
	signal NextState											: T_STATE;
	attribute FSM_ENCODING	of State			: signal is getFSMEncoding_gray(DEBUG);

	signal FISTypeRegister								: T_SATA_FISTYPE									:= SATA_FISTYPE_UNKNOWN;
	signal FlagRegister										: T_SLV_8													:= (others => '0');
	signal StatusRegister									: T_SLV_8													:= (others => '0');
	signal EndStatusRegister							: T_SLV_8													:= (others => '0');
	signal ErrorRegister									: T_SLV_8													:= (others => '0');
	signal AddressRegister								: T_SLV_48												:= (others => '0');
	signal SectorCountRegister						: T_SLV_16												:= (others => '0');
	signal TransferCountRegister					: T_SLV_16												:= (others => '0');

	signal FISTypeRegister_rst						: std_logic;
	signal FISTypeRegister_en							: std_logic;
	signal FlagRegister_en								: std_logic;
	signal StatusRegister_en							: std_logic;
	signal EndStatusRegister_en						: std_logic;
	signal ErrorRegister_en								: std_logic;
	signal AddressRegister_en0						: std_logic;
	signal AddressRegister_en8						: std_logic;
	signal AddressRegister_en16						: std_logic;
	signal AddressRegister_en24						: std_logic;
	signal AddressRegister_en32						: std_logic;
	signal AddressRegister_en40						: std_logic;
	signal SectorCountRegister_en0				: std_logic;
	signal SectorCountRegister_en8				: std_logic;
	signal TransferCountRegister_en				: std_logic;

begin

	process(Clock)
	begin
		if rising_edge(Clock) then
			if (Reset = '1') then
				State			<= ST_RESET;
			else
				State			<= NextState;
			end if;
		end if;
	end process;

	process(State, Link_Status, FISTypeRegister, Link_RX_Valid, Link_RX_Data, Link_RX_SOF, Link_RX_EOF, Link_RX_FS_Valid, Link_RX_FS_CRCOK, Link_RX_FS_SyncEsc, RX_Ack	)
	begin
		NextState										<= State;

		Status											<= SATA_FISD_STATUS_RECEIVING;

		Link_RX_Ack									<= '0';
		Link_RX_FS_Ack							<= '0';

		RX_Data											<= Link_RX_Data;
		RX_SOP											<= '0';
		RX_EOP											<= '0';
		RX_Valid										<= '0';

		FISTypeRegister_rst					<= '0';
		FISTypeRegister_en					<= '0';
		FlagRegister_en							<= '0';
		StatusRegister_en						<= '0';
		EndStatusRegister_en				<= '0';
		ErrorRegister_en						<= '0';
		AddressRegister_en0					<= '0';
		AddressRegister_en8					<= '0';
		AddressRegister_en16				<= '0';
		AddressRegister_en24				<= '0';
		AddressRegister_en32				<= '0';
		AddressRegister_en40				<= '0';
		SectorCountRegister_en0			<= '0';
		SectorCountRegister_en8			<= '0';
		TransferCountRegister_en		<= '0';

		UpdateATARegisters					<= '0';

		case State is
			when ST_RESET =>
				-- Clock might be unstable is this state. In this case either
				-- a) Reset is asserted because inital reset of the SATAController is
				--    not finished yet.
				-- b) Phy_Status is constant and not equal to SATA_LINK_STATUS_IDLE
				--    This may happen during reconfiguration due to speed negotiation.
        Status													<= SATA_FISD_STATUS_RESET;
        FISTypeRegister_rst							<= '1';

        if (Link_Status = SATA_LINK_STATUS_IDLE) then
					NextState											<= ST_IDLE;
        end if;

			when ST_IDLE =>
				Status													<= SATA_FISD_STATUS_IDLE;

				if (Link_RX_FS_Valid = '0') then
					-- wait for frame state
					null;
				elsif (Link_RX_FS_CRCOK = '1') then
					-- frame is OK and now processed
					-- wait for data frame, it's slower than frame state
					if (Link_RX_Valid = '1') then
						FISTypeRegister_en						<= '1';
						Link_RX_FS_Ack 								<= '1';
						NextState											<= ST_CHECK_FISTYPE;
					end if;
				elsif (Link_RX_FS_SyncEsc = '1') then
					Link_RX_FS_Ack 								<= '1';
					NextState											<= ST_STATUS_ERROR;
				else
					Link_RX_FS_Ack 								<= '1';
					NextState											<= ST_STATUS_CRC_ERROR;
				end if;

			when ST_CHECK_FISTYPE =>
				-- assert(Link_RX_Valid = '1')
				Status													<= SATA_FISD_STATUS_RECEIVING;

				if (Link_RX_SOF = '1') then
					Link_RX_Ack										<= '1';

					if (FISTypeRegister = SATA_FISTYPE_PIO_SETUP) then
						FlagRegister_en						<= '1';
						StatusRegister_en					<= '1';
						ErrorRegister_en					<= '1';

						if (Link_RX_EOF = '0') then
							NextState 							<= ST_FIS_PIO_SETUP_WORD_1;
						else
							NextState								<= ST_STATUS_ERROR;
						end if;

					elsif (FISTypeRegister = SATA_FISTYPE_REG_DEV_HOST) then
						FlagRegister_en						<= '1';
						StatusRegister_en					<= '1';
						ErrorRegister_en					<= '1';

						if (Link_RX_EOF = '0') then
							NextState 							<= ST_FIS_REG_DEV_HOST_WORD_1;
						else
							NextState								<= ST_STATUS_ERROR;
						end if;

					elsif (FISTypeRegister = SATA_FISTYPE_DMA_ACTIVATE) then
						if (Link_RX_EOF = '1') then
							NextState 							<= ST_RECEIVE_OK;
						else
							NextState 							<= ST_DISCARD_FRAME_1;
						end if;

					elsif (FISTypeRegister = SATA_FISTYPE_DATA) then
						if (Link_RX_EOF = '0') then
							NextState 							<= ST_FIS_DATA_1;						-- goto Data FIS processing
						else
							NextState								<= ST_STATUS_ERROR;
						end if;
					else
						if (Link_RX_EOF = '0') then
							NextState								<= ST_DISCARD_FRAME_1;
						else
							NextState								<= ST_STATUS_ERROR;
						end if;
					end if;	-- FISType_i
				else	-- Link_RX_SOF
					NextState										<= ST_DISCARD_FRAME_1;
				end if;

			-- ============================================================
			-- register transfer: device => host
			-- ============================================================
			when ST_FIS_REG_DEV_HOST_WORD_1 =>
				if (Link_RX_Valid = '1') then
					Link_RX_Ack										<= '1';

					AddressRegister_en0						<= '1';
					AddressRegister_en16					<= '1';
					AddressRegister_en32					<= '1';
					-- DeviceNumber / Heads

					if (Link_RX_EOF = '0') then
						NextState 									<= ST_FIS_REG_DEV_HOST_WORD_2;
					else
						NextState										<= ST_STATUS_ERROR;
					end if;
				end if;

			when ST_FIS_REG_DEV_HOST_WORD_2 =>
				if (Link_RX_Valid = '1') then
					Link_RX_Ack										<= '1';

					AddressRegister_en8						<= '1';
					AddressRegister_en24					<= '1';
					AddressRegister_en40					<= '1';

					if (Link_RX_EOF = '0') then
						NextState 									<= ST_FIS_REG_DEV_HOST_WORD_3;
					else
						NextState										<= ST_STATUS_ERROR;
					end if;
				end if;

			when ST_FIS_REG_DEV_HOST_WORD_3 =>
				if (Link_RX_Valid = '1') then
					Link_RX_Ack										<= '1';

					SectorCountRegister_en0				<= '1';
					SectorCountRegister_en8				<= '1';

					if (Link_RX_EOF = '0') then
						NextState 									<= ST_FIS_REG_DEV_HOST_WORD_4;
					else
						NextState										<= ST_STATUS_ERROR;
					end if;
				end if;

			when ST_FIS_REG_DEV_HOST_WORD_4 =>
				if (Link_RX_Valid = '1') then
					Link_RX_Ack										<= '1';

					if (Link_RX_EOF = '1') then
						UpdateATARegisters					<= '1';
						NextState 									<= ST_RECEIVE_OK;
					else
						NextState										<= ST_STATUS_ERROR;
					end if;
				end if;

			-- ============================================================
			-- PIO Setup
			-- ============================================================
			when ST_FIS_PIO_SETUP_WORD_1 =>
				if (Link_RX_Valid = '1') then
					Link_RX_Ack										<= '1';

					AddressRegister_en0						<= '1';
					AddressRegister_en16					<= '1';
					AddressRegister_en32					<= '1';
					-- DeviceNumber / Heads

					if (Link_RX_EOF = '0') then
						NextState 									<= ST_FIS_PIO_SETUP_WORD_2;
					else
						NextState										<= ST_STATUS_ERROR;
					end if;
				end if;

			when ST_FIS_PIO_SETUP_WORD_2 =>
				if (Link_RX_Valid = '1') then
					Link_RX_Ack										<= '1';

					AddressRegister_en8						<= '1';
					AddressRegister_en24					<= '1';
					AddressRegister_en40					<= '1';

					if (Link_RX_EOF = '0') then
						NextState 									<= ST_FIS_PIO_SETUP_WORD_3;
					else
						NextState										<= ST_STATUS_ERROR;
					end if;
				end if;

			when ST_FIS_PIO_SETUP_WORD_3 =>
				if (Link_RX_Valid = '1') then
					Link_RX_Ack										<= '1';

					SectorCountRegister_en0				<= '1';
					SectorCountRegister_en8				<= '1';
					EndStatusRegister_en					<= '1';

					if (Link_RX_EOF = '0') then
						NextState 									<= ST_FIS_PIO_SETUP_WORD_4;
					else
						NextState										<= ST_STATUS_ERROR;
					end if;
				end if;

			when ST_FIS_PIO_SETUP_WORD_4 =>
				if (Link_RX_Valid = '1') then
					Link_RX_Ack										<= '1';

					TransferCountRegister_en			<= '1';

					if (Link_RX_EOF = '1') then
						UpdateATARegisters					<= '1';
						NextState 									<= ST_RECEIVE_OK;
					else
						NextState 									<= ST_DISCARD_FRAME_1;
					end if;
				end if;

			-- ============================================================
			-- Data
			-- ============================================================
			when ST_FIS_DATA_1 =>
				-- passthrought handshaking signals
				RX_Valid												<= Link_RX_Valid;
				Link_RX_Ack											<= RX_Ack;
        RX_EOP                          <= Link_RX_EOF;
				RX_SOP													<= '1';

				-- if streaming is possible => stream first Word; set SOP; goto DATA_N
				if ((Link_RX_Valid = '1') and (RX_Ack = '1')) then
					if (Link_RX_EOF = '1') then
						NextState 									<= ST_RECEIVE_OK;
					else	-- EOF
						NextState										<= ST_FIS_DATA_N;
					end if;
				end if;

			when ST_FIS_DATA_N =>
				RX_Valid												<= Link_RX_Valid;
				Link_RX_Ack											<= RX_Ack;
        RX_EOP                          <= Link_RX_EOF;

				-- if streaming is possible => stream first Word; set SOP; goto DATA_N
				if ((Link_RX_Valid = '1') and (RX_Ack = '1')) then
					if (Link_RX_EOF = '1') then
						NextState 									<= ST_RECEIVE_OK;
					end if;
				end if;

			when ST_RECEIVE_OK =>
				Status													<= SATA_FISD_STATUS_RECEIVE_OK;
				FISTypeRegister_rst							<= '1';
				NextState												<= ST_IDLE;

			when ST_STATUS_ERROR =>
				Status													<= SATA_FISD_STATUS_ERROR;
				FISTypeRegister_rst							<= '1';
				NextState												<= ST_IDLE;

			when ST_STATUS_CRC_ERROR =>
				Status													<= SATA_FISD_STATUS_CRC_ERROR;
				FISTypeRegister_rst							<= '1';
				NextState												<= ST_IDLE;


			-- ============================================================
			-- Discard remaining frame
			-- ============================================================
			when ST_DISCARD_FRAME_1 =>
				Status													<= SATA_FISD_STATUS_ERROR;
				Link_RX_Ack											<= '1';

				if ((Link_RX_Valid = '1') and (Link_RX_EOF = '1')) then
					FISTypeRegister_rst						<= '1';
					NextState 										<= ST_IDLE;
				else
					NextState											<= ST_DISCARD_FRAME_N;
				end if;

			when ST_DISCARD_FRAME_N =>
				Status													<= SATA_FISD_STATUS_DISCARD_FRAME;
				Link_RX_Ack											<= '1';

				if ((Link_RX_Valid = '1') and (Link_RX_EOF = '1')) then
					FISTypeRegister_rst						<= '1';
					NextState 										<= ST_IDLE;
				end if;

		end case;
	end process;

	-- ================================================================
	-- ATA registers - temporary saved
	-- ================================================================
	process(Clock)
	begin
		if rising_edge(Clock) then
			if (FISTypeRegister_rst = '1') then
				FISTypeRegister	<= SATA_FISTYPE_UNKNOWN;
			elsif (FISTypeRegister_en = '1') then
				FISTypeRegister	<= to_sata_fistype(Alias_FISType);
			end if;

			-- FlagRegister
			if (FlagRegister_en	= '1') then
				FlagRegister		<= Alias_FlagReg;
			end if;

			-- StatusRegister
			if (StatusRegister_en	= '1') then
				StatusRegister	<= Alias_StatusReg;
			end if;

			-- EndStatusRegister
			if (EndStatusRegister_en	= '1') then
				EndStatusRegister	<= Alias_EndStatusReg;
			end if;

			-- ErrorRegister
			if (ErrorRegister_en	= '1') then
				ErrorRegister	<= Alias_ErrorReg;
			end if;

			-- AddressRegister
			if (AddressRegister_en0	= '1') then
				AddressRegister(7 downto 0)	<= Alias_LBA0;
			end if;

			if (AddressRegister_en8	= '1') then
				AddressRegister(15 downto 8)	<= Alias_LBA8;
			end if;

			if (AddressRegister_en16	= '1') then
				AddressRegister(23 downto 16)	<= Alias_LBA16;
			end if;

			if (AddressRegister_en24	= '1') then
				AddressRegister(31 downto 24)	<= Alias_LBA24;
			end if;

			if (AddressRegister_en32	= '1') then
				AddressRegister(39 downto 32)	<= Alias_LBA32;
			end if;

			if (AddressRegister_en40	= '1') then
				AddressRegister(47 downto 40)	<= Alias_LBA40;
			end if;

			-- SectorCountRegister
			if (SectorCountRegister_en0	= '1') then
				SectorCountRegister(7 downto 0)		<= Alias_SecCount0;
			end if;

			if (SectorCountRegister_en8	= '1') then
				SectorCountRegister(15 downto 8)	<= Alias_SecCount8;
			end if;

			-- TransferCountRegister
			if (TransferCountRegister_en	= '1') then
				TransferCountRegister				<= Alias_TransferCount;
			end if;
		end if;
	end process;

	FISType															<= FISTypeRegister;

	ATADeviceRegisters.Flags						<= to_sata_ata_device_flags(FlagRegister);
	ATADeviceRegisters.Status						<= to_sata_ata_device_register_status(StatusRegister);
	ATADeviceRegisters.EndStatus				<= to_sata_ata_device_register_status(EndStatusRegister);
	ATADeviceRegisters.Error						<= to_sata_ata_device_register_error(ErrorRegister);
	ATADeviceRegisters.LBlockAddress		<= AddressRegister;
	ATADeviceRegisters.SectorCount			<= SectorCountRegister;
	ATADeviceRegisters.TransferCount		<= TransferCountRegister when (TransferCountRegister_en = '0') else Alias_TransferCount;

	-- debug ports
	-- ==========================================================================================================================================================
	genDebug : if (ENABLE_DEBUGPORT = TRUE) generate
		function dbg_EncodeState(st : T_STATE) return std_logic_vector is
		begin
			return to_slv(T_STATE'pos(st), log2ceilnz(T_STATE'pos(T_STATE'high) + 1));
		end function;

	begin
		genXilinx : if (VENDOR = VENDOR_XILINX) generate
			function dbg_GenerateStateEncodings return string is
				variable  l : STD.TextIO.line;
			begin
				for i in T_STATE loop
					STD.TextIO.write(l, str_replace(T_STATE'image(i), "st_", ""));
					STD.TextIO.write(l, ';');
				end loop;
				return  l.all;
			end function;

			function dbg_GenerateStatusEncodings return string is
				variable  l : STD.TextIO.line;
			begin
				for i in T_SATA_FISDECODER_STATUS loop
					STD.TextIO.write(l, str_replace(T_SATA_FISDECODER_STATUS'image(i), "sata_fisd_status_", ""));
					STD.TextIO.write(l, ';');
				end loop;
				return  l.all;
			end function;

--			constant dummy : T_BOOLVEC := (
--				0 => dbg_ExportEncoding("Transport Layer FIS-Decoder - FSM", dbg_GenerateStateEncodings,  PROJECT_DIR & "ChipScope/TokenFiles/FSM_TransLayer_FISD.tok"),
--				1 => dbg_ExportEncoding("Transport Layer FIS-Decoder - Status", dbg_GenerateStatusEncodings,  PROJECT_DIR & "ChipScope/TokenFiles/ENUM_Trans_FISD_Status.tok")
--			);
		begin
		end generate;

		DebugPortOut.FSM		<= dbg_EncodeState(State);
	end generate;
end;
