library IEEE;
use			IEEE.STD_LOGIC_1164.all;
use			IEEE.NUMERIC_STD.all;

library PoC;
use			PoC.config.all;
use			PoC.utils.all;

library L_Global;
use			PoC.GlobalTypes.all;

package EthDebug is


end;

package body EthDebug is

end package body;