LIBRARY IEEE;
USE			IEEE.STD_LOGIC_1164.ALL;
USE			IEEE.NUMERIC_STD.ALL;

LIBRARY PoC;
USE			PoC.functions.ALL;

LIBRARY	L_Global;
USE			L_Global.GlobalTypes.ALL;

-- Usage
-- ====================================
-- LIBRARY L_SATAController;
-- USE L_SATAController.SATATypes.ALL;

PACKAGE SATATypes IS
	-- declare attributes
	ATTRIBUTE ENUM_ENCODING	: STRING;
	

-- ==================================================================
-- link layer types
-- ==================================================================
	TYPE T_SATA_LINK_COMMAND IS (
		SATA_LINK_CMD_NONE,
		SATA_LINK_CMD_RESET
	);

	TYPE T_SATA_LINK_STATUS IS (
		SATA_LINK_STATUS_IDLE,
		SATA_LINK_STATUS_SENDING,
		SATA_LINK_STATUS_RECEIVING,
		SATA_LINK_STATUS_COMMUNICATION_ERROR,
		SATA_LINK_STATUS_ERROR
	);
	
	TYPE T_SATA_LINK_ERROR IS (
		SATA_LINK_ERROR_NONE,
		SATA_LINK_ERROR_PHY_COMRESET,
		SATA_LINK_ERROR_PHY_8B10B_ERROR,
		SATA_LINK_ERROR_LINK_RXFIFO_FULL,
		SATA_LINK_ERROR_LINK_FSM
	);
	
	TYPE T_SATA_PRIMITIVE IS (					-- Primitive Name				Byte 3,	Byte 2,	Byte 1,	Byte 0
		SATA_PRIMITIVE_NONE,							-- no primitive
		SATA_PRIMITIVE_ALIGN,							-- ALIGN								D27.3,	D10.2,	D10.2,	K28.5
		SATA_PRIMITIVE_SYNC,							-- SYNC									D21.5,	D21.5,	D21.4,	K28.3
		SATA_PRIMITIVE_DIAL_TONE,					-- D10.2								D10.2,	D10.2,	D10.2,	D10.2
		SATA_PRIMITIVE_SOF,								-- SOF									D23.1,	D23.1,	D21.5,	K28.3
		SATA_PRIMITIVE_EOF,								-- EOF									D21.6,	D21.6,	D21.5,	K28.3
		SATA_PRIMITIVE_HOLD,							-- HOLD									D21.6,	D21.6,	D10.5,	K28.3
		SATA_PRIMITIVE_HOLD_ACK,					-- HOLDA								D21.4,	D21.4,	D10.5,	K28.3
		SATA_PRIMITIVE_CONT,							-- CONT									D25.4,	D25.4,	D10.5,	K28.3
		SATA_PRIMITIVE_R_OK,							-- R_OK									D21.1,	D21.1,	D21.5,	K28.3
		SATA_PRIMITIVE_R_ERROR,						-- R_ERR								D22.2,	D22.2,	D21.5,	K28.3
		SATA_PRIMITIVE_R_IP,							-- R_IP									D21.2,	D21.2,	D21.5,	K28.3
		SATA_PRIMITIVE_RX_RDY,						-- R_RDY								D10.2,	D10.2,	D21.4,	K28.3
		SATA_PRIMITIVE_TX_RDY,						-- X_RDY								D23.2,	D23.2,	D21.5,	K28.3
		SATA_PRIMITIVE_DMA_TERM,					-- DMAT									D22.1,	D22.1,	D21.5,	K28.3
		SATA_PRIMITIVE_WAIT_TERM,					-- WTRM									D24.2,	D24.2,	D21.5,	K28.3
		SATA_PRIMITIVE_PM_ACK,						-- PMACK								D
		SATA_PRIMITIVE_PM_NACK,						-- PMNAK								D
		SATA_PRIMITIVE_PM_REQ_P,					-- PMREQ_P							D	
		SATA_PRIMITIVE_PM_REQ_S,					-- PMREQ_S							D	
		SATA_PRIMITIVE_ILLEGAL
	);
	CONSTANT T_SATA_PRIMITIVE_COUNT		: INTEGER										:= T_SATA_PRIMITIVE'pos(SATA_PRIMITIVE_ILLEGAL) + 1;

	CONSTANT SATA_MAX_FRAMESIZE_B			: POSITIVE									:= 8192;
	CONSTANT SATA_WORD_BW							: POSITIVE									:= 32;

	TYPE T_SATA_LINK_COMMAND_VECTOR		IS ARRAY (NATURAL RANGE <>) OF T_SATA_LINK_COMMAND;
	TYPE T_SATA_LINK_STATUS_VECTOR		IS ARRAY (NATURAL RANGE <>) OF T_SATA_LINK_STATUS;
	TYPE T_SATA_LINK_ERROR_VECTOR			IS ARRAY (NATURAL RANGE <>) OF T_SATA_LINK_ERROR;

-- ==================================================================
-- physical layer types
-- ==================================================================
	SUBTYPE T_SATA_GENERATION				IS INTEGER RANGE 0 TO 5;
	
	CONSTANT SATA_GENERATION_1			: T_SATA_GENERATION		:= 0;
	CONSTANT SATA_GENERATION_2			: T_SATA_GENERATION		:= 1;
	CONSTANT SATA_GENERATION_3			: T_SATA_GENERATION		:= 2;
	CONSTANT SATA_GENERATION_AUTO		: T_SATA_GENERATION		:= 4;
	CONSTANT SATA_GENERATION_ERROR	: T_SATA_GENERATION		:= 5;
	
--	ATTRIBUTE ENUM_ENCODING OF T_SATA_GENERATION	: TYPE IS "00 01 10 11";
	
	TYPE T_SATA_PHY_COMMAND IS (
		SATA_PHY_CMD_NONE,					-- no command
		SATA_PHY_CMD_RESET,					-- reset retry and generation counter => reprogramm to initial configuration
		SATA_PHY_CMD_NEWLINK_UP			-- reset retry counter use same generation
	);

	TYPE T_SATA_PHY_STATUS IS (
		SATA_PHY_STATUS_RESET,
		SATA_PHY_STATUS_LINK_UP,
		SATA_PHY_STATUS_LINK_OK,
		SATA_PHY_STATUS_LINK_BROKEN,
		SATA_PHY_STATUS_RECEIVED_RESET,
		SATA_PHY_STATUS_CHANGE_SPEED,
		SATA_PHY_STATUS_ERROR							-- FIXME: unused?
	);

	-- FIXME: unused?
	TYPE T_SATA_PHY_ERROR IS (
		SATA_PHY_ERROR_NONE,
		SATA_PHY_ERROR_COMRESET,
		SATA_PHY_ERROR_LINK_DEAD,
		SATA_PHY_ERROR_NEGOTIATION_ERROR,
		SATA_PHY_ERROR_FSM
	);

	TYPE T_SGEN_SGEN								IS ARRAY (T_SATA_GENERATION) OF T_SATA_GENERATION;			-- REFACTOR:
	TYPE T_SGEN2_SGEN								IS ARRAY (T_SATA_GENERATION) OF T_SGEN_SGEN;						-- REFACTOR:
	TYPE T_SGEN3_SGEN								IS ARRAY (T_SATA_GENERATION) OF T_SGEN2_SGEN;						-- REFACTOR:
	
	TYPE T_SGEN_INT									IS ARRAY (T_SATA_GENERATION) OF INTEGER;								-- REFACTOR:
	TYPE T_SGEN2_INT								IS ARRAY (T_SATA_GENERATION) OF T_SGEN_INT;							-- REFACTOR:
	
	TYPE T_SATA_GENERATION_VECTOR		IS ARRAY (NATURAL RANGE <>) OF T_SATA_GENERATION;
	TYPE T_SATA_PHY_COMMAND_VECTOR	IS ARRAY (NATURAL RANGE <>) OF T_SATA_PHY_COMMAND;
	TYPE T_SATA_PHY_STATUS_VECTOR		IS ARRAY (NATURAL RANGE <>) OF T_SATA_PHY_STATUS;
	TYPE T_SATA_PHY_ERROR_VECTOR		IS ARRAY (NATURAL RANGE <>) OF T_SATA_PHY_ERROR;


-- ==================================================================
-- transceiver types
-- ==================================================================
	-- oob signals
	TYPE T_SATA_OOB IS (
		SATA_OOB_NONE,
		SATA_OOB_READY,
		SATA_OOB_COMRESET,
		SATA_OOB_COMWAKE
	);
	
	-- CharIsK
	SUBTYPE T_SATA_CIK2		IS STD_LOGIC_VECTOR(1 DOWNTO 0);			-- REFACTOR: to v5 gtp
	SUBTYPE T_SATA_CIK		IS STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	-- transceiver commands
	TYPE T_SATA_TRANSCEIVER_COMMAND IS (
		SATA_TRANSCEIVER_CMD_NONE,
		SATA_TRANSCEIVER_CMD_POWERDOWN,
		SATA_TRANSCEIVER_CMD_POWERUP,
		SATA_TRANSCEIVER_CMD_RESET,
		SATA_TRANSCEIVER_CMD_RECONFIG,
		SATA_TRANSCEIVER_CMD_UNLOCK
	);
	
	-- transceiver status
	TYPE T_SATA_TRANSCEIVER_STATUS IS (
		SATA_TRANSCEIVER_STATUS_POWERED_DOWN,
		SATA_TRANSCEIVER_STATUS_RESETING,
		SATA_TRANSCEIVER_STATUS_RECONFIGURING,
		SATA_TRANSCEIVER_STATUS_RELOADING,
		SATA_TRANSCEIVER_STATUS_READY,
		SATA_TRANSCEIVER_STATUS_READY_LOCKED,
		SATA_TRANSCEIVER_STATUS_NO_DEVICE,
		SATA_TRANSCEIVER_STATUS_NEW_DEVICE,
		SATA_TRANSCEIVER_STATUS_ERROR
	);

	-- transceiver error
	TYPE T_SATA_TRANSCEIVER_ERROR IS (
		SATA_TRANSCEIVER_ERROR_NONE,
		SATA_TRANSCEIVER_ERROR_FSM
	);

	-- transmitter errors
	TYPE T_SATA_TRANSCEIVER_TX_ERROR IS (
		SATA_TRANSCEIVER_TX_ERROR_NONE,
		SATA_TRANSCEIVER_TX_ERROR_ENCODER,
		SATA_TRANSCEIVER_TX_ERROR_BUFFER
	);
	
	-- receiver errors
	TYPE T_SATA_TRANSCEIVER_RX_ERROR IS (
		SATA_TRANSCEIVER_RX_ERROR_NONE,
		SATA_TRANSCEIVER_RX_ERROR_ALIGNEMENT,
		SATA_TRANSCEIVER_RX_ERROR_DISPARITY,
		SATA_TRANSCEIVER_RX_ERROR_DECODER,
		SATA_TRANSCEIVER_RX_ERROR_BUFFER
	);

	TYPE T_SATA_CIK2_VECTOR										IS ARRAY (NATURAL RANGE <>) OF T_SATA_CIK2;			-- REFACTOR: to v5 gtp
	TYPE T_SATA_CIK_VECTOR										IS ARRAY (NATURAL RANGE <>) OF T_SATA_CIK;
	TYPE T_SATA_OOB_VECTOR										IS ARRAY (NATURAL RANGE <>) OF T_SATA_OOB;
	TYPE T_SATA_TRANSCEIVER_COMMAND_VECTOR		IS ARRAY (NATURAL RANGE <>) OF T_SATA_TRANSCEIVER_COMMAND;
	TYPE T_SATA_TRANSCEIVER_STATUS_VECTOR			IS ARRAY (NATURAL RANGE <>) OF T_SATA_TRANSCEIVER_STATUS;
	TYPE T_SATA_TRANSCEIVER_TX_ERROR_VECTOR		IS ARRAY (NATURAL RANGE <>) OF T_SATA_TRANSCEIVER_TX_ERROR;
	TYPE T_SATA_TRANSCEIVER_RX_ERROR_VECTOR		IS ARRAY (NATURAL RANGE <>) OF T_SATA_TRANSCEIVER_RX_ERROR;

-- ==================================================================
--common sata types
-- ==================================================================
	TYPE T_SATA_COMMAND IS (
		SATA_CMD_NONE,
		SATA_CMD_RESET,
		SATA_CMD_RESET_CONNECTION,				-- invoke COMRESET / COMINIT
		SATA_CMD_RESET_LINKLAYER,					-- reset LinkLayer => send SYNC-primitive
		SATA_CMD_POWERDOWN
	);

	TYPE T_SATA_STATUS IS RECORD
		LinkLayer							: T_SATA_LINK_STATUS;
		PhysicalLayer					: T_SATA_PHY_STATUS;
		TransceiverLayer			: T_SATA_TRANSCEIVER_STATUS;
	END RECORD;
	
	TYPE T_SATA_ERROR IS RECORD
		LinkLayer							: T_SATA_LINK_ERROR;
		PhysicalLayer					: T_SATA_PHY_ERROR;
		TransceiverLayer_TX		: T_SATA_TRANSCEIVER_TX_ERROR;
		TransceiverLayer_RX		: T_SATA_TRANSCEIVER_RX_ERROR;
	END RECORD;

	TYPE T_SATA_DEVICE_TYPE IS (
		SATA_DEVICE_TYPE_HOST,
		SATA_DEVICE_TYPE_DEVICE
	);
	
	TYPE T_SATA_COMMAND_VECTOR				IS ARRAY (NATURAL RANGE <>) OF  T_SATA_COMMAND;
	TYPE T_SATA_STATUS_VECTOR					IS ARRAY (NATURAL RANGE <>) OF  T_SATA_STATUS;
	TYPE T_SATA_ERROR_VECTOR					IS ARRAY (NATURAL RANGE <>) OF  T_SATA_ERROR;
	TYPE T_SATA_DEVICE_TYPE_VECTOR		IS ARRAY (NATURAL RANGE <>) OF  T_SATA_DEVICE_TYPE;

	FUNCTION to_slv(Primitive : T_SATA_PRIMITIVE) RETURN T_SLV_32;
	
END SATATypes;


PACKAGE BODY SATATypes IS
	FUNCTION to_slv(Primitive : T_SATA_PRIMITIVE) RETURN T_SLV_32 IS
	BEGIN																														--																							K symbol
																																	-- primitive name				Byte 3	Byte 2	Byte 1	Byte 0
		CASE Primitive IS																							-- =======================================================
			WHEN SATA_PRIMITIVE_NONE =>				RETURN x"00000000";				-- no primitive					
			WHEN SATA_PRIMITIVE_ALIGN =>			RETURN x"7B4A4ABC";				-- ALIGN								D27.3,	D10.2,	D10.2,	K28.5
			WHEN SATA_PRIMITIVE_SYNC =>				RETURN x"B5B5957C";				-- SYNC									D21.5,	D21.5,	D21.4,	K28.3
			WHEN SATA_PRIMITIVE_SOF =>				RETURN x"3737B57C";				-- SOF									D23.1,	D23.1,	D21.5,	K28.3
			WHEN SATA_PRIMITIVE_EOF =>				RETURN x"D5D5B57C";				-- EOF									D21.6,	D21.6,	D21.5,	K28.3
			WHEN SATA_PRIMITIVE_HOLD =>				RETURN x"D5D5AA7C";				-- HOLD									D21.6,	D21.6,	D10.5,	K28.3
			WHEN SATA_PRIMITIVE_HOLD_ACK =>		RETURN x"9595AA7C";				-- HOLDA								D21.4,	D21.4,	D10.5,	K28.3
			WHEN SATA_PRIMITIVE_CONT =>				RETURN x"9999AA7C";				-- CONT									D25.4,	D25.4,	D10.5,	K28.3
			WHEN SATA_PRIMITIVE_R_OK =>				RETURN x"3535B57C";				-- R_OK									D21.1,	D21.1,	D21.5,	K28.3
			WHEN SATA_PRIMITIVE_R_ERROR =>		RETURN x"5656B57C";				-- R_ERR								D22.2,	D22.2,	D21.5,	K28.3
			WHEN SATA_PRIMITIVE_R_IP =>				RETURN x"5555B57C";				-- R_IP									D21.2,	D21.2,	D21.5,	K28.3
			WHEN SATA_PRIMITIVE_RX_RDY =>			RETURN x"4A4A957C";				-- R_RDY								D10.2,	D10.2,	D21.4,	K28.3
			WHEN SATA_PRIMITIVE_TX_RDY =>			RETURN x"5757B57C";				-- X_RDY								D23.2,	D23.2,	D21.5,	K28.3
			WHEN SATA_PRIMITIVE_DMA_TERM =>		RETURN x"3636B57C";				-- DMAT									D22.1,	D22.1,	D21.5,	K28.3
			WHEN SATA_PRIMITIVE_WAIT_TERM =>	RETURN x"5858B57C";				-- WTRM									D24.2,	D24.2,	D21.5,	K28.3
			WHEN SATA_PRIMITIVE_PM_ACK =>			RETURN x"9595957C";				-- PMACK								D21.4,	D21.4,	D21.4,	K28.3
			WHEN SATA_PRIMITIVE_PM_NACK =>		RETURN x"F5F5957C";				-- PMNAK								D21.7,	D21.7,	D21.4,	K28.3
			WHEN SATA_PRIMITIVE_PM_REQ_P =>		RETURN x"1717B57C";				-- PMREQ_P							D23.0,	D23.0,	D21.5,	K28.3
			WHEN SATA_PRIMITIVE_PM_REQ_S =>		RETURN x"7575957C";				-- PMREQ_S							D21.3,	D21.3,	D21.4,	K28.3
			WHEN SATA_PRIMITIVE_DIAL_TONE =>	RETURN x"4A4A4A4A";				-- 											D10.2,	D10.2,	D10.2,	D10.2
			WHEN SATA_PRIMITIVE_ILLEGAL =>		RETURN (OTHERS => 'X');		-- "ERROR"
		END CASE;
	END;
	
END PACKAGE BODY;
