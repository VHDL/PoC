-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- =============================================================================
-- Authors:         Stefan Unrein
--
-- Entity:          A generic AXI4-Lite version register for Git.
--
-- Description:
-- -------------------------------------
-- This version register can be auto filled with constants from Git. Software
-- can read from what revision a firmware (bitstream, PL code) was build.
--
-- Use the pre-synthesis script from
--     PoC/tools/git/preSynth_GitVersionRegister_Vivado.tcl
-- to create a memory file with all necessary information. Add this file name to
-- the VERSION_FILE_NAME generic.
--
-- License:
-- =============================================================================
-- Copyright 2024-2025 The PoC-Library Authors
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--    http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- =============================================================================

library IEEE;
use     IEEE.std_logic_1164.all;
use     IEEE.numeric_std.all;

use     work.config.all;
use     work.utils.all;
use     work.vectors.all;
use     work.strings.all;
use     work.axi4lite.all;
use     work.xil.all;

use     work.mem_GitVersionRegister.all;


entity AXI4Lite_GitVersionRegister is
	Generic (
		VERSION_FILE_NAME     : string;                                                      -- Path to version-memory generated by preSynth_GitVersionRegister_Vivado.tcl
		WRITE_FILE_NAME       : string  := "";                                               -- Writes the Version-Register structure to a csv file with this name. Leave empty if not used.
		INCLUDE_XIL_DNA       : boolean := false;                                            -- Enable Xilinx DNA Port
		INCLUDE_XIL_USER_EFUSE : boolean := false;                                            -- Enable Xilinx User eFuse
		USER_ID               : std_logic_vector(95 downto 0) := (others => '0');            -- User ID saved in register "UID.User_ID"
		IGNORE_HIGH_ADDRESS               : boolean         := true;                         -- Disables the High-Address Check. If the Base-Address of the whole register can be ignored, leave as true, otherwhise, the addresses in the config need be set with base-address
		RESPONSE_ON_ERROR                 : T_AXI4_Response := C_AXI4_RESPONSE_DECODE_ERROR  -- If not address matches then config of the AXI4Lite transaction, return this code
	);
	Port (
		Clock        : in  std_logic;
		Reset        : in  std_logic;

		AXI4Lite_m2s : in  T_AXI4Lite_BUS_M2S;
		AXI4Lite_s2m : out T_AXI4Lite_BUS_S2M
	);
end entity;


architecture rtl of AXI4Lite_GitVersionRegister is
	constant CONFIG      : T_AXI4_Register_Vector       := get_Version_Descriptor;
	constant VersionData : T_SLVV_32(0 to C_Num_Version_Header - 1) := read_Version_from_mem(PROJECT_DIR & VERSION_FILE_NAME);

	signal   RegisterFile_ReadPort   : T_SLVV(0 to CONFIG'Length -1)(DATA_BITS - 1 downto 0);
	signal   RegisterFile_WritePort  : T_SLVV(0 to CONFIG'Length -1)(DATA_BITS - 1 downto 0);

	signal   UID_vec                 : T_SLVV(0 to C_Num_Reg_UID -1)(DATA_BITS - 1 downto 0);

begin
	Header_file_gen : if WRITE_FILE_NAME'length > 0 generate
	begin
		assert write_csv_file(PROJECT_DIR & WRITE_FILE_NAME, CONFIG) report "Failure in writing CSV File" severity warning;
	end generate;

	AXI4LiteReg : entity work.AXI4Lite_Register
	generic map(
		CONFIG                  => CONFIG,
		IGNORE_HIGH_ADDRESS     => IGNORE_HIGH_ADDRESS,
		RESPONSE_ON_ERROR       => RESPONSE_ON_ERROR
	)
	port map(
		Clock                   => Clock,
		Reset                   => Reset,

		AXI4Lite_m2s            => AXI4Lite_m2s,
		AXI4Lite_s2m            => AXI4Lite_s2m,

		RegisterFile_ReadPort   => RegisterFile_ReadPort,
		RegisterFile_WritePort  => RegisterFile_WritePort
	);
	RegisterFile_WritePort(0 to C_Num_Version_Header -1) <= VersionData;
	RegisterFile_WritePort(C_Num_Version_Header to C_Num_Version_Register -1) <= UID_vec;

	---------------------------------
	-- Generate data for UID-vector
	---------------------------------
	UID_vec(low(C_Num_reg_UID_vec, 2) to high(C_Num_reg_UID_vec, 2)) <= to_slvv_32(USER_ID);

	dna_gen : if INCLUDE_XIL_DNA generate
		signal DNA : std_logic_vector(get_DNABITS -1 downto 0);
	begin
		DNA_inst : component xil_DNAPort
		port map(
			Clock   => Clock,
			Reset   => Reset,
			Valid   => open,
			DataOut => DNA
		);
		UID_vec(low(C_Num_reg_UID_vec, 0) to high(C_Num_reg_UID_vec, 0)) <= rev(to_slvv_32(resize(DNA, C_Num_reg_UID_vec(0) * 32)));
	else generate
		UID_vec(low(C_Num_reg_UID_vec, 0) to high(C_Num_reg_UID_vec, 0)) <= (others => (others => '0'));
	end generate;

	efuse_gen : if INCLUDE_XIL_USER_EFUSE generate
		assert false report "AXI4Lite_GitVersionRegister:: INCLUDE_XIL_USR_EFUSE is currently not supported, feel free to implement it ;)" severity failure;
	else generate
		UID_vec(low(C_Num_reg_UID_vec, 1) to high(C_Num_reg_UID_vec, 1)) <= (others => (others => '0'));
	end generate;
end architecture;
