-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- 
-- ============================================================================
-- Package:					Project specific configuration.
-- 
-- Authors:         Thomas B. Preusser
--                  Martin Zabel
--                  Patrick Lehmann
--
-- Description:
-- ------------------------------------
--		This is a template file. 
--		The global package common/config evaluates the settings declared in this file.
--
-- Usage:
--		1) Copy this file into your project's source directory and rename it to my_config.vhdl.
--		2) Add file to library "poc" in your synthesis tool.
--		3) Change setup appropriately.
--
-- License:
-- ============================================================================
-- Copyright 2007-2014 Technische Universitaet Dresden - Germany
--										 Chair for VLSI-Design, Diagnostics and Architecture
-- 
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
-- 
--    http://www.apache.org/licenses/LICENSE-2.0
-- 
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- ============================================================================

library PoC;

package my_config is
  -- Change these lines to setup configuration.
  constant MY_BOARD		: string := "ML605";								-- ML605 - Xilinx Virtex 6 reference design board: XC6VLX240T
  constant MY_DEVICE	: string := "None";									-- infer from MY_BOARD
 
end my_config;

package body my_config is

end my_config;