-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- 
-- =============================================================================
-- Package:					TODO
--
-- Authors:					Patrick Lehmann
--
-- Description:
-- ------------------------------------
--		TODO
-- 
-- License:
-- =============================================================================
-- Copyright 2007-2014 Technische Universitaet Dresden - Germany
--										 Chair for VLSI-Design, Diagnostics and Architecture
-- 
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
-- 
--		http://www.apache.org/licenses/LICENSE-2.0
-- 
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- =============================================================================

LIBRARY IEEE;
USE			IEEE.STD_LOGIC_1164.ALL;
USE			IEEE.NUMERIC_STD.ALL;

LIBRARY PoC;
USE			PoC.utils.ALL;
USE			PoC.vectors.ALL;
--USE			PoC.strings.ALL;
--USE			PoC.sata.ALL;


ENTITY sata_CommandFSM IS
	GENERIC (
		DEBUG															: BOOLEAN								:= FALSE;
		SIM_EXECUTE_IDENTIFY_DEVICE				: BOOLEAN								:= TRUE				-- required by CommandLayer: load device parameters
	);
	PORT (
		Clock															: IN	STD_LOGIC;
		Reset															: IN	STD_LOGIC;

		-- for measurement purposes only
		Config_BurstSize									: IN	T_SLV_16;

		-- ATAStreamingController interface
		Command														: IN	T_ATA_CMD_COMMAND;
		Status														: OUT	T_ATA_CMD_STATUS;
		Error															: OUT	T_ATA_CMD_ERROR;

		Address_LB												: IN	T_SLV_48;
		BlockCount_LB											: IN	T_SLV_48;

		TX_en															: OUT	STD_LOGIC;

		RX_SOR														: OUT	STD_LOGIC;
		RX_EOR														: OUT	STD_LOGIC;

		-- TransporTrans interface
		Trans_Command											: OUT	T_SATA_TRANS_COMMAND;
		Trans_Status											: IN	T_SATA_TRANS_STATUS;
		Trans_Error												: IN	T_SATA_TRANS_ERROR;
		
		Trans_UpdateATAHostRegisters			: OUT STD_LOGIC;
		Trans_ATAHostRegisters						: OUT T_ATA_HOST_REGISTERS;
		
		Trans_RX_SOT											: IN	STD_LOGIC;
		Trans_RX_EOT											: IN	STD_LOGIC;
		
		-- IdentifyDeviceFilter interface
		IDF_Enable												: OUT	STD_LOGIC;
		IDF_DriveInformation							: IN	T_DRIVE_INFORMATION;
		IDF_Error													: IN	STD_LOGIC
	);
END;

ARCHITECTURE rtl OF sata_CommandFSM IS
	ATTRIBUTE KEEP												: BOOLEAN;
	ATTRIBUTE FSM_ENCODING								: STRING;

	CONSTANT MAX_BLOCKCOUNT								: POSITIVE												:= ite(SIMULATION, SIM_MAX_BLOCKCOUNT, ATA_MAX_BLOCKCOUNT);

	-- 1 => single transfer
	-- F => first transfer
	-- N => next transfer
	-- L => last transfer
	TYPE T_STATE IS (
		ST_RESET,
		ST_INIT,
		ST_IDLE,
		ST_IDENTIFY_DEVICE_WAIT,	ST_IDENTIFY_DEVICE_CHECK,
		ST_READ_1_WAIT,		ST_READ_F_WAIT,		ST_READ_N_WAIT,		ST_READ_L_WAIT,
		ST_WRITE_1_WAIT,	ST_WRITE_F_WAIT,	ST_WRITE_N_WAIT,	ST_WRITE_L_WAIT,
		ST_FLUSH_CACHE_WAIT,
		ST_ERROR
	);
	
	SIGNAL State													: T_STATE													:= ST_RESET;
	SIGNAL NextState											: T_STATE;
	ATTRIBUTE FSM_ENCODING	OF State			: SIGNAL IS ite(DEBUG					, "gray", ite((VENDOR = VENDOR_XILINX), "auto", "default"));
	
	SIGNAL Trans_Command_i								: T_SATA_TRANS_COMMAND;
	
	SIGNAL Load														: STD_LOGIC;
	SIGNAL NextTransfer										: STD_LOGIC;
	SIGNAL LastTransfer										: STD_LOGIC;
	SIGNAL BurstCount_us									: UNSIGNED(16 DOWNTO 0);
	SIGNAL Address_LB_us									: UNSIGNED(47 DOWNTO 0);
	SIGNAL Address_LB_us_d								: UNSIGNED(47 DOWNTO 0)						:= (OTHERS => '0');
	SIGNAL Address_LB_us_d_nx							: UNSIGNED(47 DOWNTO 0);
	SIGNAL BlockCount_LB_us								: UNSIGNED(47 DOWNTO 0);
	SIGNAL BlockCount_LB_us_d							: UNSIGNED(47 DOWNTO 0)						:= (OTHERS => '0');
	SIGNAL BlockCount_LB_us_d_nx					: UNSIGNED(47 DOWNTO 0);
	
	SIGNAL ATA_Address_LB_us							: UNSIGNED(47 DOWNTO 0);
	SIGNAL ATA_BlockCount_LB_us						: UNSIGNED(15 DOWNTO 0);
	
	SIGNAL ATA_Address_LB									: T_SLV_48;
	SIGNAL ATA_BlockCount_LB							: T_SLV_16;
	
	ATTRIBUTE KEEP OF Load								: SIGNAL IS DEBUG					;
	ATTRIBUTE KEEP OF NextTransfer				: SIGNAL IS DEBUG					;
	ATTRIBUTE KEEP OF LastTransfer				: SIGNAL IS DEBUG					;
	
BEGIN
-- ATA_Device_register => TD=0 -> 40   / TD=1 -> 50

	PROCESS(Clock)
	BEGIN
		IF rising_edge(Clock) THEN
			IF (Reset = '1') THEN
				State			<= ST_RESET;
			ELSE
				State			<= NextState;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS(State, Command, Trans_Status, IDF_Error, IDF_DriveInformation, ATA_Address_LB, ATA_BlockCount_LB, LastTransfer, Trans_RX_SOT, Trans_RX_EOT)
	BEGIN
		NextState																		<= State;
		
		Status																			<= ATA_CMD_STATUS_RESET; -- just in case
		Error																				<= ATA_CMD_ERROR_NONE;
		
		Load																				<= '0';
		NextTransfer																<= '0';
		
		TX_en																				<= '0';
		
		RX_SOR																			<= '0';
		RX_EOR																			<= '0';
		
		Trans_Command_i															<= SATA_TRANS_CMD_NONE;
		Trans_UpdateATAHostRegisters								<= '0';
		Trans_ATAHostRegisters.Flag_C								<= '0';
		Trans_ATAHostRegisters.Command							<= to_slv(ATA_CMD_NONE);			-- Command register
		Trans_ATAHostRegisters.Control							<= (OTHERS => '0');						-- Control register
		Trans_ATAHostRegisters.Feature							<= (OTHERS => '0');						-- Feature register
		Trans_ATAHostRegisters.LBlockAddress				<= (OTHERS => '0');						-- logical block address (LBA)
		Trans_ATAHostRegisters.SectorCount					<= (OTHERS => '0');						-- 
		
		IDF_Enable																	<= '0';
		
		CASE State IS
			WHEN ST_RESET =>
				Status																			<= ATA_CMD_STATUS_RESET;
        
        IF (Trans_Status = SATA_TRANS_STATUS_IDLE) THEN
					IF (SIM_EXECUTE_IDENTIFY_DEVICE = TRUE) THEN
						NextState																<= ST_INIT;
					ELSE
						NextState																<= ST_IDLE;
					END IF;
        END IF;
			
			WHEN ST_INIT =>
        -- assert Trans_Status = SATA_TRANS_STATUS_IDLE
				Status																			<= ATA_CMD_STATUS_INITIALIZING;
						
				-- TransferLayer
				Trans_Command_i															<= SATA_TRANS_CMD_TRANSFER;
				Trans_UpdateATAHostRegisters								<= '1';
				Trans_ATAHostRegisters.Flag_C								<= '1';
				Trans_ATAHostRegisters.Command							<= to_slv(ATA_CMD_IDENTIFY_DEVICE);			-- Command register
				Trans_ATAHostRegisters.Control							<= (OTHERS => '0');											-- Control register
				Trans_ATAHostRegisters.Feature							<= (OTHERS => '0');											-- Feature register
				Trans_ATAHostRegisters.LBlockAddress				<= (OTHERS => '0');											-- logical block address (LBA)
				Trans_ATAHostRegisters.SectorCount					<= (OTHERS => '0');											-- 
			
				-- IdentifyDeviceFilter
				IDF_Enable																	<= '1';
			
				NextState																		<= ST_IDENTIFY_DEVICE_WAIT;
			
			WHEN ST_IDLE =>
        -- assert Trans_Status = SATA_TRANS_STATUS_IDLE
				Status																			<= ATA_CMD_STATUS_IDLE;
			
				CASE Command IS
					WHEN ATA_CMD_CMD_NONE =>
						NULL;
						
					WHEN ATA_CMD_CMD_RESET =>
						NULL;
					
					WHEN ATA_CMD_CMD_IDENTIFY_DEVICE =>
						Status																	<= ATA_CMD_STATUS_EXECUTING;
						
						-- TransferLayer
						Trans_Command_i													<= SATA_TRANS_CMD_TRANSFER;
						Trans_UpdateATAHostRegisters						<= '1';
						Trans_ATAHostRegisters.Flag_C						<= '1';
						Trans_ATAHostRegisters.Command					<= to_slv(ATA_CMD_IDENTIFY_DEVICE);			-- Command register
						Trans_ATAHostRegisters.Control					<= (OTHERS => '0');											-- Control register
						Trans_ATAHostRegisters.Feature					<= (OTHERS => '0');											-- Feature register
						Trans_ATAHostRegisters.LBlockAddress		<= (OTHERS => '0');											-- logical block address (LBA)
						Trans_ATAHostRegisters.SectorCount			<= (OTHERS => '0');											-- 
					
						-- IdentifyDeviceFilter
						IDF_Enable															<= '1';
					
						NextState																<= ST_IDENTIFY_DEVICE_WAIT;
						
					WHEN ATA_CMD_CMD_READ =>
						Status																	<= ATA_CMD_STATUS_RECEIVING;
		
						-- TransferGenerator
						Load																		<= '1';
						
						-- TransferLayer
						Trans_Command_i													<= SATA_TRANS_CMD_TRANSFER;
						Trans_UpdateATAHostRegisters						<= '1';
						Trans_ATAHostRegisters.Flag_C						<= '1';
						Trans_ATAHostRegisters.Command					<= to_slv(ATA_CMD_DMA_READ_EXT);				-- Command register
						Trans_ATAHostRegisters.Control					<= (OTHERS => '0');											-- Control register
						Trans_ATAHostRegisters.Feature					<= (OTHERS => '0');											-- Feature register
						Trans_ATAHostRegisters.LBlockAddress		<= ATA_Address_LB;											-- logical block address (LBA)
						Trans_ATAHostRegisters.SectorCount			<= ATA_BlockCount_LB;										-- 
			
						IF (LastTransfer = '0') THEN
							NextState															<= ST_READ_F_WAIT;
						ELSE
							NextState															<= ST_READ_1_WAIT;
						END IF;
						
					WHEN ATA_CMD_CMD_WRITE =>
						Status																	<= ATA_CMD_STATUS_SENDING;
						
						-- TransferGenerator
						Load																		<= '1';
						
						-- TransferLayer
						Trans_Command_i													<= SATA_TRANS_CMD_TRANSFER;
						Trans_UpdateATAHostRegisters						<= '1';
						Trans_ATAHostRegisters.Flag_C						<= '1';
						Trans_ATAHostRegisters.Command					<= to_slv(ATA_CMD_DMA_WRITE_EXT);				-- Command register
						Trans_ATAHostRegisters.Control					<= (OTHERS => '0');											-- Control register
						Trans_ATAHostRegisters.Feature					<= (OTHERS => '0');											-- Feature register
						Trans_ATAHostRegisters.LBlockAddress		<= ATA_Address_LB;											-- logical block address (LBA)
						Trans_ATAHostRegisters.SectorCount			<= ATA_BlockCount_LB;										-- 
			
						IF (LastTransfer = '0') THEN
							NextState															<= ST_WRITE_F_WAIT;
						ELSE
							NextState															<= ST_WRITE_1_WAIT;
						END IF;

					WHEN ATA_CMD_CMD_FLUSH_CACHE =>
						IF (IDF_DriveInformation.Valid = '0') THEN
							Status																<= ATA_CMD_STATUS_INITIALIZING;
						ELSE
							Status																<= ATA_CMD_STATUS_EXECUTING;
						END IF;
						
						-- TransferLayer
						Trans_Command_i													<= SATA_TRANS_CMD_TRANSFER;
						Trans_UpdateATAHostRegisters						<= '1';
						Trans_ATAHostRegisters.Flag_C						<= '1';
						Trans_ATAHostRegisters.Command					<= to_slv(ATA_CMD_FLUSH_CACHE_EXT);			-- Command register
						Trans_ATAHostRegisters.Control					<= (OTHERS => '0');											-- Control register
						Trans_ATAHostRegisters.Feature					<= (OTHERS => '0');											-- Feature register
						Trans_ATAHostRegisters.LBlockAddress		<= (OTHERS => '0');											-- logical block address (LBA)
						Trans_ATAHostRegisters.SectorCount			<= (OTHERS => '0');											-- 
			
						NextState																<= ST_FLUSH_CACHE_WAIT;
						
					WHEN OTHERS =>
						Status																	<= ATA_CMD_STATUS_ERROR;
						Error																		<= ATA_CMD_ERROR_FSM;
						NextState																<= ST_ERROR;

				END CASE;
			
			WHEN ST_IDENTIFY_DEVICE_WAIT =>
				IF (IDF_DriveInformation.Valid = '0') THEN
					Status																		<= ATA_CMD_STATUS_INITIALIZING;
				ELSE
					Status																		<= ATA_CMD_STATUS_EXECUTING;
				END IF;
			
				IDF_Enable																	<= '1';
				
				IF (Trans_Status = SATA_TRANS_STATUS_TRANSFERING) THEN
					IF (IDF_Error = '1') THEN
						Status																	<= ATA_CMD_STATUS_ERROR;
						Error																		<= ATA_CMD_ERROR_IDENTIFY_DEVICE_ERROR;
						NextState																<= ST_ERROR;
					END IF;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_TRANSFER_OK) THEN
					IF (IDF_Error = '0') THEN
						NextState																<= ST_IDENTIFY_DEVICE_CHECK;
					ELSE
						Status																	<= ATA_CMD_STATUS_ERROR;
						Error																		<= ATA_CMD_ERROR_IDENTIFY_DEVICE_ERROR;
						NextState																<= ST_ERROR;
					END IF;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_ERROR) THEN
					Status																		<= ATA_CMD_STATUS_ERROR;
					Error																			<= ATA_CMD_ERROR_TRANSPORT_ERROR;
					NextState																	<= ST_ERROR;
				END IF;
				
			WHEN ST_IDENTIFY_DEVICE_CHECK =>
				Status																			<= ATA_CMD_STATUS_INITIALIZING;
			
				IF (IDF_DriveInformation.Valid = '1') THEN
					IF ((IDF_DriveInformation.ATACapabilityFlags.SupportsDMA = '1') AND
							(IDF_DriveInformation.ATACapabilityFlags.SupportsLBA = '1') AND
							(IDF_DriveInformation.ATACapabilityFlags.Supports48BitLBA = '1') AND
							(IDF_DriveInformation.ATACapabilityFlags.SupportsFLUSH_CACHE = '1') AND
							(IDF_DriveInformation.ATACapabilityFlags.SupportsFLUSH_CACHE_EXT = '1')) THEN
						NextState																<= ST_IDLE;
					ELSE	-- device not supported
						Status																	<= ATA_CMD_STATUS_ERROR;
						Error																		<= ATA_CMD_ERROR_DEVICE_NOT_SUPPORTED;
						NextState																<= ST_ERROR;
					END IF;
				ELSE
					-- information are not valid
					Status																		<= ATA_CMD_STATUS_ERROR;
					Error																			<= ATA_CMD_ERROR_IDENTIFY_DEVICE_ERROR;
					NextState																	<= ST_ERROR;
				END IF;
				
			-- ============================================================
			-- ATA command: ATA_CMD_CMD_READ
			-- ============================================================
			WHEN ST_READ_1_WAIT =>
				Status																	<= ATA_CMD_STATUS_RECEIVING;
				
				RX_SOR																	<= Trans_RX_SOT;
				RX_EOR																	<= Trans_RX_EOT;
				
				IF (Trans_Status = SATA_TRANS_STATUS_TRANSFERING) THEN
					NULL;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_TRANSFER_OK) THEN
					NextState															<= ST_IDLE;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_ERROR) THEN
					Status																<= ATA_CMD_STATUS_ERROR;
					Error																	<= ATA_CMD_ERROR_TRANSPORT_ERROR;
					NextState															<= ST_ERROR;
				END IF;
			
			WHEN ST_READ_F_WAIT =>
				Status																	<= ATA_CMD_STATUS_RECEIVING;
				
				RX_SOR																	<= Trans_RX_SOT;
				
				IF (Trans_Status = SATA_TRANS_STATUS_TRANSFERING) THEN
					NULL;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_TRANSFER_OK) THEN
					-- TransferGenerator
					NextTransfer													<= '1';
					
					-- TransferLayer
					Trans_Command_i												<= SATA_TRANS_CMD_TRANSFER;
					Trans_UpdateATAHostRegisters					<= '1';
					Trans_ATAHostRegisters.Flag_C					<= '1';
					Trans_ATAHostRegisters.Command				<= to_slv(ATA_CMD_DMA_READ_EXT);				-- Command register
					Trans_ATAHostRegisters.Control				<= (OTHERS => '0');											-- Control register
					Trans_ATAHostRegisters.Feature				<= (OTHERS => '0');											-- Feature register
					Trans_ATAHostRegisters.LBlockAddress	<= ATA_Address_LB;											-- logical block address (LBA)
					Trans_ATAHostRegisters.SectorCount		<= ATA_BlockCount_LB;										-- 
					
					IF (LastTransfer = '0') THEN
						NextState														<= ST_READ_N_WAIT;
					ELSE
						NextState														<= ST_READ_L_WAIT;
					END IF;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_ERROR) THEN
					Status																<= ATA_CMD_STATUS_ERROR;
					Error																	<= ATA_CMD_ERROR_TRANSPORT_ERROR;
					NextState															<= ST_ERROR;
				END IF;
			
			WHEN ST_READ_N_WAIT =>
				Status																	<= ATA_CMD_STATUS_RECEIVING;
				
				IF (Trans_Status = SATA_TRANS_STATUS_TRANSFERING) THEN
					NULL;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_TRANSFER_OK) THEN
					-- TransferGenerator
					NextTransfer													<= '1';
					
					-- TransferLayer
					Trans_Command_i												<= SATA_TRANS_CMD_TRANSFER;
					Trans_UpdateATAHostRegisters					<= '1';
					Trans_ATAHostRegisters.Flag_C					<= '1';
					Trans_ATAHostRegisters.Command				<= to_slv(ATA_CMD_DMA_READ_EXT);				-- Command register
					Trans_ATAHostRegisters.Control				<= (OTHERS => '0');											-- Control register
					Trans_ATAHostRegisters.Feature				<= (OTHERS => '0');											-- Feature register
					Trans_ATAHostRegisters.LBlockAddress	<= ATA_Address_LB;											-- logical block address (LBA)
					Trans_ATAHostRegisters.SectorCount		<= ATA_BlockCount_LB;										-- 
					
					IF (LastTransfer = '0') THEN
						NextState														<= ST_READ_N_WAIT;
					ELSE
						NextState														<= ST_READ_L_WAIT;
					END IF;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_ERROR) THEN
					Status																<= ATA_CMD_STATUS_ERROR;
					Error																	<= ATA_CMD_ERROR_TRANSPORT_ERROR;
					NextState															<= ST_ERROR;
				END IF;
			
			WHEN ST_READ_L_WAIT =>
				Status																	<= ATA_CMD_STATUS_RECEIVING;
				
				RX_EOR																	<= Trans_RX_EOT;
				
				IF (Trans_Status = SATA_TRANS_STATUS_TRANSFERING) THEN
					NULL;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_TRANSFER_OK) THEN
					NextState															<= ST_IDLE;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_ERROR) THEN
					Status																<= ATA_CMD_STATUS_ERROR;
					Error																	<= ATA_CMD_ERROR_TRANSPORT_ERROR;
					NextState															<= ST_ERROR;
				END IF;
			
			-- ============================================================
			-- ATA command: ATA_CMD_CMD_WRITE
			-- ============================================================
			WHEN ST_WRITE_1_WAIT =>
				Status																	<= ATA_CMD_STATUS_SENDING;
				TX_en																		<= '1';
				
				IF (Trans_Status = SATA_TRANS_STATUS_TRANSFERING) THEN
					NULL;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_TRANSFER_OK) THEN
					NextState															<= ST_IDLE;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_ERROR) THEN
					Status																<= ATA_CMD_STATUS_ERROR;
					Error																	<= ATA_CMD_ERROR_TRANSPORT_ERROR;
					NextState															<= ST_ERROR;
				END IF;
				
			WHEN ST_WRITE_F_WAIT =>
				Status																	<= ATA_CMD_STATUS_SENDING;
				TX_en																		<= '1';
				
				IF (Trans_Status = SATA_TRANS_STATUS_TRANSFERING) THEN
					NULL;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_TRANSFER_OK) THEN
					-- TransferGenerator
					NextTransfer													<= '1';
					
					-- TransferLayer
					Trans_Command_i												<= SATA_TRANS_CMD_TRANSFER;
					Trans_UpdateATAHostRegisters					<= '1';
					Trans_ATAHostRegisters.Flag_C					<= '1';
					Trans_ATAHostRegisters.Command				<= to_slv(ATA_CMD_DMA_WRITE_EXT);				-- Command register
					Trans_ATAHostRegisters.Control				<= (OTHERS => '0');											-- Control register
					Trans_ATAHostRegisters.Feature				<= (OTHERS => '0');											-- Feature register
					Trans_ATAHostRegisters.LBlockAddress	<= ATA_Address_LB;											-- logical block address (LBA)
					Trans_ATAHostRegisters.SectorCount		<= ATA_BlockCount_LB;										-- 
					
					IF (LastTransfer = '0') THEN
						NextState														<= ST_WRITE_N_WAIT;
					ELSE
						NextState														<= ST_WRITE_L_WAIT;
					END IF;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_ERROR) THEN
					Status																<= ATA_CMD_STATUS_ERROR;
					Error																	<= ATA_CMD_ERROR_TRANSPORT_ERROR;
					NextState															<= ST_ERROR;
				END IF;
			
			WHEN ST_WRITE_N_WAIT =>
				Status																	<= ATA_CMD_STATUS_SENDING;
				TX_en																		<= '1';
				
				IF (Trans_Status = SATA_TRANS_STATUS_TRANSFERING) THEN
					NULL;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_TRANSFER_OK) THEN
					-- TransferGenerator
					NextTransfer													<= '1';
					
					-- TransferLayer
					Trans_Command_i												<= SATA_TRANS_CMD_TRANSFER;
					Trans_UpdateATAHostRegisters					<= '1';
					Trans_ATAHostRegisters.Flag_C					<= '1';
					Trans_ATAHostRegisters.Command				<= to_slv(ATA_CMD_DMA_WRITE_EXT);				-- Command register
					Trans_ATAHostRegisters.Control				<= (OTHERS => '0');											-- Control register
					Trans_ATAHostRegisters.Feature				<= (OTHERS => '0');											-- Feature register
					Trans_ATAHostRegisters.LBlockAddress	<= ATA_Address_LB;											-- logical block address (LBA)
					Trans_ATAHostRegisters.SectorCount		<= ATA_BlockCount_LB;										-- 
					
					IF (LastTransfer = '0') THEN
						NextState														<= ST_WRITE_N_WAIT;
					ELSE
						NextState														<= ST_WRITE_L_WAIT;
					END IF;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_ERROR) THEN
					Status																<= ATA_CMD_STATUS_ERROR;
					Error																	<= ATA_CMD_ERROR_TRANSPORT_ERROR;
					NextState															<= ST_ERROR;
				END IF;
			
			WHEN ST_WRITE_L_WAIT =>
				Status																	<= ATA_CMD_STATUS_SENDING;
				TX_en																		<= '1';
				
				IF (Trans_Status = SATA_TRANS_STATUS_TRANSFERING) THEN
					NULL;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_TRANSFER_OK) THEN
					NextState															<= ST_IDLE;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_ERROR) THEN
					Status																<= ATA_CMD_STATUS_ERROR;
					Error																	<= ATA_CMD_ERROR_TRANSPORT_ERROR;
					NextState															<= ST_ERROR;
				END IF;
		
			-- ============================================================
			-- ATA command: ATA_CMD_CMD_FLUSH_CACHE
			-- ============================================================
			WHEN ST_FLUSH_CACHE_WAIT =>
				Status																	<= ATA_CMD_STATUS_EXECUTING;
				
				IF (Trans_Status = SATA_TRANS_STATUS_TRANSFERING) THEN
					NULL;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_TRANSFER_OK) THEN
					NextState															<= ST_IDLE;
				ELSIF (Trans_Status = SATA_TRANS_STATUS_ERROR) THEN
					Status																<= ATA_CMD_STATUS_ERROR;
					Error																	<= ATA_CMD_ERROR_TRANSPORT_ERROR;
					NextState															<= ST_ERROR;
				END IF;

			WHEN ST_ERROR =>
				Status																	<= ATA_CMD_STATUS_ERROR;
				Error																		<= ATA_CMD_ERROR_FSM;

		END CASE;
	END PROCESS;
	
	Trans_Command				<= Trans_Command_i WHEN rising_edge(Clock);
	
	-- transfer and address generation
	Address_LB_us				<= unsigned(Address_LB);
	BlockCount_LB_us		<= unsigned(BlockCount_LB);
	
	LastTransfer				<= to_sl(ite((Load = '1'), BlockCount_LB_us, BlockCount_LB_us_d) <= BurstCount_us);
	
	PROCESS(Load, LastTransfer, Address_LB_us, BlockCount_LB_us, Address_LB_us_d, BlockCount_LB_us_d, Address_LB_us_d_nx, BlockCount_LB_us_d_nx, Config_BurstSize)
	BEGIN
		IF (Load = '1') THEN
			Address_LB_us_d_nx														<= Address_LB_us;
			BlockCount_LB_us_d_nx													<= BlockCount_LB_us;
		ELSE
			Address_LB_us_d_nx														<= Address_LB_us_d;
			BlockCount_LB_us_d_nx													<= BlockCount_LB_us_d;
		END IF;

		ATA_Address_LB_us			<= Address_LB_us_d_nx;
		
		IF (LastTransfer = '0') THEN
			IF (MAX_BLOCKCOUNT = unsigned(Config_BurstSize)) THEN
				ATA_BlockCount_LB_us												<= (OTHERS => '0');
			ELSE
				ATA_BlockCount_LB_us												<= unsigned(Config_BurstSize);													-- => ATA_MAX_BLOCKCOUNT is encoded as 0x0000000000
			END IF;
		ELSE
			ATA_BlockCount_LB_us													<= BlockCount_LB_us_d_nx(ATA_BlockCount_LB_us'range);		--
		END IF;
	END PROCESS;

	ATA_Address_LB				<= std_logic_vector(ATA_Address_LB_us);
	ATA_BlockCount_LB			<= std_logic_vector(ATA_BlockCount_LB_us);
	
	BurstCount_us					<= ite((Config_BurstSize = (Config_BurstSize'range => '0')), to_unsigned(MAX_BLOCKCOUNT, BurstCount_us'length), unsigned('0' & Config_BurstSize));
	
	PROCESS(Clock)
	BEGIN
		IF rising_edge(Clock) THEN
			IF (Reset = '1') THEN
				Address_LB_us_d						<= (OTHERS => '0');
				BlockCount_LB_us_d				<= (OTHERS => '0');
			ELSE
				IF ((Load = '1') OR (NextTransfer = '1')) THEN
					Address_LB_us_d					<= Address_LB_us_d_nx			+ BurstCount_us;
					BlockCount_LB_us_d			<= BlockCount_LB_us_d_nx	- BurstCount_us;
				END IF;
			END IF;
		END IF;
	END PROCESS;
END;
