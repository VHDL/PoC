-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- 
-- ============================================================================
-- Package:					This VHDL package declares new physical types and their
--									conversion functions.
--
-- Authors:					Patrick Lehmann
-- 
-- Description:
-- ------------------------------------
--		For detailed documentation see below.
--	
--		NAMING CONVENTION:
--			t - time
--			p - period
--			d - delay
--			f - frequency
--			br - baud rate
--			vec - vector
--			
--		ATTENTION:
--			This package is not supported by Xilinx Synthese Tools prior to 14.x!
--			
--			It was successfully tested with:
--				- Xilinx Synthesis Tool (XST) 14.7 and Xilinx ISE Simulator (iSim) 14.7
--				- Xilinx Vivado	Synthesis 2014.2 and Xilinx Vivado Simulator (xSim) 2014.2
--				- Quartus II 13.1
--				- QuestaSim 10.0d
--				- GHDL 0.31
--		
-- License:
-- ============================================================================
-- Copyright 2007-2014 Technische Universitaet Dresden - Germany,
--										 Chair for VLSI-Design, Diagnostics and Architecture
-- 
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
-- 
--		http://www.apache.org/licenses/LICENSE-2.0
-- 
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- ============================================================================

library PoC;
use			PoC.my_config.MY_VERBOSE;
use			PoC.strings.all;


package physical is
	
	type FREQ is range 0 to INTEGER'high units
		Hz;
		kHz = 1000 Hz;
		MHz = 1000 kHz;
		GHz = 1000 MHz;
		THz = 1000 GHz;
	end units;

	type BAUD is range 0 to INTEGER'high units
		Bd;
		kBd = 1000 Bd;
		MBd = 1000 kBd;
		GBd = 1000 MBd;
	end units;

	type MEMORY is range 0 to INTEGER'high units
		B;
		KiB = 1000 B;
		MiB = 1000 KiB;
		GiB = 1000 MiB;
		TiB = 1000 GiB;
	end units;
	
	SUBTYPE	T_DELAY							IS TIME;
	SUBTYPE	T_PERIOD						IS TIME;																	-- see QUESTIONs below
	TYPE		T_TIMEVEC						IS ARRAY(NATURAL RANGE <>) OF TIME;				-- use short VEC names (see PoC.utils T_INTVEC) or long forms (like STD_LOGIC_VECTOR)?
	TYPE		T_FREQVEC						IS ARRAY(NATURAL RANGE <>) OF FREQ;
	TYPE		T_BAUDVEC						IS ARRAY(NATURAL RANGE <>) OF BAUD;
	TYPE		T_MEMVEC						IS ARRAY(NATURAL RANGE <>) OF MEMORY;
	
	function to_time(f : FREQ)	return TIME;
	function to_freq(p : TIME)	return FREQ;
	function to_freq(br : BAUD)	return FREQ;
	
	-- if-then-else
	function ite(cond : BOOLEAN; value1 : TIME;	value2 : TIME) return TIME;
	function ite(cond : BOOLEAN; value1 : FREQ;	value2 : FREQ) return FREQ;
	function ite(cond : BOOLEAN; value1 : BAUD;	value2 : BAUD) return BAUD;
	function ite(cond : BOOLEAN; value1 : MEMORY;	value2 : MEMORY) return MEMORY;
	
	-- min/ max for 2 arguments
	function min(arg1 : TIME; arg2 : TIME) return TIME;						-- Calculates: min(arg1, arg2) for times
	function min(arg1 : FREQ; arg2 : FREQ) return FREQ;						-- Calculates: min(arg1, arg2) for frequencies
	function min(arg1 : BAUD; arg2 : BAUD) return BAUD;						-- Calculates: min(arg1, arg2) for symbols per second
	function min(arg1 : MEMORY; arg2 : MEMORY) return MEMORY;			-- Calculates: min(arg1, arg2) for memory
	
	function max(arg1 : TIME; arg2 : TIME) return TIME;						-- Calculates: max(arg1, arg2) for times
	function max(arg1 : FREQ; arg2 : FREQ) return FREQ;						-- Calculates: max(arg1, arg2) for frequencies
	function max(arg1 : BAUD; arg2 : BAUD) return BAUD;						-- Calculates: max(arg1, arg2) for symbols per second
	function max(arg1 : MEMORY; arg2 : MEMORY) return MEMORY;			-- Calculates: max(arg1, arg2) for memory
	
	-- min/max/sum as vector aggregation
	function min(vec : T_TIMEVEC)	return TIME;										-- Calculates: min(vec) for a time vector
	function min(vec : T_FREQVEC)	return FREQ;										-- Calculates: min(vec) for a frequency vector
	function min(vec : T_BAUDVEC)	return BAUD;										-- Calculates: min(vec) for a baud vector
	function min(vec : T_MEMVEC)	return MEMORY;									-- Calculates: min(vec) for a memory vector
	
	function max(vec : T_TIMEVEC)	return TIME;										-- Calculates: max(vec) for a time vector
	function max(vec : T_FREQVEC)	return FREQ;										-- Calculates: max(vec) for a frequency vector
	function max(vec : T_BAUDVEC)	return BAUD;										-- Calculates: max(vec) for a baud vector
	function max(vec : T_MEMVEC)	return MEMORY;									-- Calculates: max(vec) for a memory vector
	
	-- QUESTION: some sum functions are not meaningful -> orthogonal function/type system
	function sum(vec : T_TIMEVEC)	return TIME;										-- Calculates: sum(vec) for a time vector
	function sum(vec : T_FREQVEC)	return FREQ;										-- Calculates: sum(vec) for a frequency vector
	function sum(vec : T_BAUDVEC)	return BAUD;										-- Calculates: sum(vec) for a baud vector
	function sum(vec : T_MEMVEC)	return MEMORY;									-- Calculates: sum(vec) for a memory vector
	
	-- convert standard types (NATURAL, REAL) to time (TIME)
	function fs2Time(t_fs : NATURAL)		return TIME;
	function ps2Time(t_ps : NATURAL)		return TIME;
	function ns2Time(t_ns : NATURAL)		return TIME;
	function us2Time(t_us : NATURAL)		return TIME;
	function ms2Time(t_ms : NATURAL)		return TIME;
	function sec2Time(t_sec : NATURAL)	return TIME;
	
	function fs2Time(t_fs : REAL)				return TIME;
	function ps2Time(t_ps : REAL)				return TIME;
	function ns2Time(t_ns : REAL)				return TIME;
	function us2Time(t_us : REAL)				return TIME;
	function ms2Time(t_ms : REAL)				return TIME;
	function sec2Time(t_sec : REAL)			return TIME;
	
	-- convert standard types (NATURAL, REAL) to period (TIME)
	-- QUESTION: rename 'Time' to 'Period' and change result type to 'PERIOD' (<=> subtype of TIME)
	function Hz2Time(f_Hz : NATURAL)		return TIME;
	function kHz2Time(f_kHz : NATURAL)	return TIME;
	function MHz2Time(f_MHz : NATURAL)	return TIME;
	function GHz2Time(f_GHz : NATURAL)	return TIME;
	function THz2Time(f_THz : NATURAL)	return TIME;

	function Hz2Time(f_Hz : REAL)				return TIME;
	function kHz2Time(f_kHz : REAL) 		return TIME;
	function MHz2Time(f_MHz : REAL) 		return TIME;
	function GHz2Time(f_GHz : REAL) 		return TIME;
	function THz2Time(f_THz : REAL) 		return TIME;
	
	-- convert standard types (NATURAL, REAL) to frequency (FREQ)
	function Hz2Freq(f_Hz : NATURAL)		return FREQ;
	function kHz2Freq(f_kHz : NATURAL)	return FREQ;
	function MHz2Freq(f_MHz : NATURAL)	return FREQ;
	function GHz2Freq(f_GHz : NATURAL)	return FREQ;
	function THz2Freq(f_THz : NATURAL)	return FREQ;
	
	function Hz2Freq(f_Hz : REAL)				return FREQ;
	function kHz2Freq(f_kHz : REAL)			return FREQ;
	function MHz2Freq(f_MHz : REAL)			return FREQ;
	function GHz2Freq(f_GHz : REAL)			return FREQ;
	function THz2Freq(f_THz : REAL)			return FREQ;
	
	-- convert TIME to standard type (REAL)
	function to_real_fs(t : TIME)				return REAL;
	function to_real_ps(t : TIME)				return REAL;
	function to_real_ns(t : TIME)				return REAL;
	function to_real_us(t : TIME)				return REAL;
	function to_real_ms(t : TIME)				return REAL;
	function to_real_sec(t : TIME)			return REAL;

	-- convert FREQ to standard type (REAL)
	function to_real_Hz(f : FREQ) 			return REAL;
	function to_real_kHz(f : FREQ)			return REAL;
	function to_real_MHz(f : FREQ)			return REAL;
	function to_real_GHz(f : FREQ)			return REAL;
	function to_real_THz(f : FREQ)			return REAL;

	-- convert physical types (TIME, FREQ) to standard type (REAL)
	-- QUESTION: alternative functions
	--	1. to_real(t : TIME; scale : T_TIMESCALE := ns), where T_TIMESCALE := enum(FS, PS, NS, ...) possible collision with physical unit names
	--	2. to_real(t : TIME; scale : TIME), example myReal := to_real(myTiming, 1 ns);
	-- 	++ less functions
	--	-- 2 parameters
	function to_real(t : TIME; scale : TIME)			return REAL;
	function to_real(f : FREQ; scale : FREQ)			return REAL;
	function to_real(f : BAUD; scale : BAUD)			return REAL;
	function to_real(f : MEMORY; scale : MEMORY)	return REAL;
	
	-- calculate needed counter cycles to achieve a given 1. timing/delay and 2. frequency/period
	-- QUESTION: if a type PERIOD (as subtype of TIME) is introduced, change TIME to PERIOD?
	function TimingToCycles(Timing : TIME; Clock_Period			: TIME) return NATURAL;
	function TimingToCycles(Timing : TIME; Clock_Frequency	: FREQ) return NATURAL;
	
	-- convert and format physical types to STRING
	function to_string(t : TIME; precision : NATURAL := 3)			return STRING;
	function to_string(f : FREQ; precision : NATURAL := 3)			return STRING;
	function to_string(br : BAUD; precision : NATURAL := 3)			return STRING;
	function to_string(mem : MEMORY; precision : NATURAL := 3)	return STRING;
	
end physical;


package body physical is
	function to_time(f : FREQ) return TIME is
		variable res : TIME;
	begin
		if		(f < 1.0 kHz) then res := (1.0 / real(f / 1.0  Hz)) * 1.0 sec;
		elsif (f < 1.0 MHz) then res := (1.0 / real(f / 1.0 kHz)) * 1.0 ms;
		elsif (f < 1.0 GHz) then res := (1.0 / real(f / 1.0 MHz)) * 1.0 us;
		elsif (f < 1.0 THz) then res := (1.0 / real(f / 1.0 GHz)) * 1.0 ns;
		else										 res := (1.0 / real(f / 1.0 THz)) * 1.0 ps;
		end if;

		assert not MY_VERBOSE report "to_time: f= " & to_string(f) & "  return " & to_string(res) severity note;
		return res;
	end function;

	function to_freq(p : TIME) return FREQ is
		variable res : FREQ;
	begin
		if		(p < 1.0 ps)	then res := (1.0 / real(p / 1.0 fs)) * 1.0 THz;
		elsif (p < 1.0 ns)	then res := (1.0 / real(p / 1.0 ps)) * 1.0 GHz;
		elsif (p < 1.0 us)	then res := (1.0 / real(p / 1.0 ns)) * 1.0 MHz;
		elsif (p < 1.0 ms)	then res := (1.0 / real(p / 1.0 us)) * 1.0 kHz;
		elsif (p < 1.0 sec) then res := (1.0 / real(p / 1.0 ms)) * 1.0  Hz;
		else report "to_freq: input period exceeds output frequency scale." severity failure;
		end if;

		assert not MY_VERBOSE report "to_freq: p= " & to_string(p) & "  return " & to_string(res) severity note;
		return res;
	end function;
	
	function to_freq(br : BAUD) return FREQ is
		variable res : FREQ;
	begin
		if		(br < 1.0 kBd) then res := (real(br / 1.0 Bd)) * 1.0  Hz;
		elsif	(br < 1.0 MBd) then res := (real(br / 1.0 kBd)) * 1.0 kHz;
		elsif	(br < 1.0 GBd) then res := (real(br / 1.0 MBd)) * 1.0 MHz;
		else											res := (real(br / 1.0 GBd)) * 1.0 GHz;
		end if;

		assert not MY_VERBOSE report "to_freq: br= " & to_string(br) & "  return " & to_string(res) severity note;
		return res;
	end function;
	
	-- if-then-else
	-- ===========================================================================
	function ite(cond : BOOLEAN; value1 : TIME;	value2 : TIME) return TIME is
	begin
		if cond then
			return value1;
		else
			return value2;
		end if;
	end function;
	
	function ite(cond : BOOLEAN; value1 : FREQ;	value2 : FREQ) return FREQ is
	begin
		if cond then
			return value1;
		else
			return value2;
		end if;
	end function;
	
	function ite(cond : BOOLEAN; value1 : BAUD;	value2 : BAUD) return BAUD is
	begin
		if cond then
			return value1;
		else
			return value2;
		end if;
	end function;
	
	function ite(cond : BOOLEAN; value1 : MEMORY;	value2 : MEMORY) return MEMORY is
	begin
		if cond then
			return value1;
		else
			return value2;
		end if;
	end function;
	
	-- min/ max for 2 arguments
	-- ===========================================================================
	-- Calculates: min(arg1, arg2) for times
	function min(arg1 : TIME; arg2 : TIME) return TIME is
	begin
		if arg1 < arg2 then return arg1; end if;
		return arg2;
	end function;
	
	-- Calculates: min(arg1, arg2) for frequencies
	function min(arg1 : FREQ; arg2 : FREQ) return FREQ is
	begin
		if arg1 < arg2 then return arg1; end if;
		return arg2;
	end function;
	
	-- Calculates: min(arg1, arg2) for symbols per second
	function min(arg1 : BAUD; arg2 : BAUD) return BAUD is
	begin
		if arg1 < arg2 then return arg1; end if;
		return arg2;
	end function;
	
	-- Calculates: min(arg1, arg2) for memory
	function min(arg1 : MEMORY; arg2 : MEMORY) return MEMORY is
	begin
		if arg1 < arg2 then return arg1; end if;
		return arg2;
	end function;
	
	-- Calculates: max(arg1, arg2) for times
	function max(arg1 : TIME; arg2 : TIME) return TIME is
	begin
		if arg1 > arg2 then return arg1; end if;
		return arg2;
	end function;

	-- Calculates: max(arg1, arg2) for frequencies
	function max(arg1 : FREQ; arg2 : FREQ) return FREQ is
	begin
		if arg1 > arg2 then return arg1; end if;
		return arg2;
	end function;

	-- Calculates: max(arg1, arg2) for symbols per second
	function max(arg1 : BAUD; arg2 : BAUD) return BAUD is
	begin
		if arg1 > arg2 then return arg1; end if;
		return arg2;
	end function;

	-- Calculates: max(arg1, arg2) for memory
	function max(arg1 : MEMORY; arg2 : MEMORY) return MEMORY is
	begin
		if arg1 > arg2 then return arg1; end if;
		return arg2;
	end function;
	
	-- min/max/sum as vector aggregation
	-- ===========================================================================
	-- Calculates: min(vec) for a time vector
	function min(vec : T_TIMEVEC)	return TIME is
		variable  res : TIME := TIME'high;
	begin
		for i in vec'range loop
			if vec(i) < res then
				res := vec(i);
			end if;
		end loop;
		return  res;
	end;
	
	-- Calculates: min(vec) for a frequency vector
	function min(vec : T_FREQVEC)	return FREQ is
		variable  res : FREQ := FREQ'high;
	begin
		for i in vec'range loop
			if vec(i) < res then
				res := vec(i);
			end if;
		end loop;
		return  res;
	end;
	
	-- Calculates: min(vec) for a baud vector
	function min(vec : T_BAUDVEC)	return BAUD is
		variable  res : BAUD := BAUD'high;
	begin
		for i in vec'range loop
			if vec(i) < res then
				res := vec(i);
			end if;
		end loop;
		return  res;
	end;
	
	-- Calculates: min(vec) for a memory vector
	function min(vec : T_MEMVEC)	return MEMORY is
		variable  res : MEMORY := MEMORY'high;
	begin
		for i in vec'range loop
			if vec(i) < res then
				res := vec(i);
			end if;
		end loop;
		return  res;
	end;
	
	-- Calculates: max(vec) for a time vector
	function max(vec : T_TIMEVEC)	return TIME is
		variable  res : TIME := TIME'low;
	begin
		for i in vec'range loop
			if vec(i) > res then
				res := vec(i);
			end if;
		end loop;
		return  res;
	end;
	
	-- Calculates: max(vec) for a frequency vector
	function max(vec : T_FREQVEC)	return FREQ is
		variable  res : FREQ := FREQ'low;
	begin
		for i in vec'range loop
			if vec(i) > res then
				res := vec(i);
			end if;
		end loop;
		return  res;
	end;
	
	-- Calculates: max(vec) for a baud vector
	function max(vec : T_BAUDVEC)	return BAUD is
		variable  res : BAUD := BAUD'low;
	begin
		for i in vec'range loop
			if vec(i) > res then
				res := vec(i);
			end if;
		end loop;
		return  res;
	end;
	
	-- Calculates: max(vec) for a memory vector
	function max(vec : T_MEMVEC)	return MEMORY is
		variable  res : MEMORY := MEMORY'low;
	begin
		for i in vec'range loop
			if vec(i) > res then
				res := vec(i);
			end if;
		end loop;
		return  res;
	end;
	
	-- Calculates: sum(vec) for a time vector
	function sum(vec : T_TIMEVEC)	return TIME is
		variable  res : TIME := 0.0 fs;
	begin
		for i in vec'range loop
			res	:= res + vec(i);
		end loop;
		return  res;
	end;
	
	-- Calculates: sum(vec) for a frequency vector
	function sum(vec : T_FREQVEC)	return FREQ is
		variable  res : FREQ := 0.0 Hz;
	begin
		for i in vec'range loop
			res	:= res + vec(i);
		end loop;
		return  res;
	end;
	
	-- Calculates: sum(vec) for a baud vector
	function sum(vec : T_BAUDVEC)	return BAUD is
		variable  res : BAUD := 0.0 Bd;
	begin
		for i in vec'range loop
			res	:= res + vec(i);
		end loop;
		return  res;
	end;
	
	-- Calculates: sum(vec) for a memory vector
	function sum(vec : T_MEMVEC)	return MEMORY is
		variable  res : MEMORY := 0.0 B;
	begin
		for i in vec'range loop
			res	:= res + vec(i);
		end loop;
		return  res;
	end;
	
	-- convert standard types (NATURAL, REAL) to time (TIME)
	-- ===========================================================================
	function fs2Time(t_fs : NATURAL) return TIME is
	begin
		return real(t_fs) * 1.0 fs;
	end function;
	
	function ps2Time(t_ps : NATURAL) return TIME is
	begin
		return real(t_ps) * 1.0 ps;
	end function;
	
	function ns2Time(t_ns : NATURAL) return TIME is
	begin
		return real(t_ns) * 1.0 ns;
	end function;
	
	function us2Time(t_us : NATURAL) return TIME is
	begin
		return real(t_us) * 1.0 us;
	end function;
	
	function ms2Time(t_ms : NATURAL) return TIME is
	begin
		return real(t_ms) * 1.0 ms;
	end function;
	
	function sec2Time(t_sec : NATURAL) return TIME is
	begin
		return real(t_sec) * 1.0 sec;
	end function;
	
	function fs2Time(t_fs : REAL) return TIME is
	begin
		return t_fs * 1.0 fs;
	end function;
	
	function ps2Time(t_ps : REAL) return TIME is
	begin
		return t_ps * 1.0 ps;
	end function;
	
	function ns2Time(t_ns : REAL) return TIME is
	begin
		return t_ns * 1.0 ns;
	end function;
	
	function us2Time(t_us : REAL) return TIME is
	begin
		return t_us * 1.0 us;
	end function;
	
	function ms2Time(t_ms : REAL) return TIME is
	begin
		return t_ms * 1.0 ms;
	end function;
	
	function sec2Time(t_sec : REAL) return TIME is
	begin
		return t_sec * 1.0 sec;
	end function;
	
	-- convert standard types (NATURAL, REAL) to period (TIME)
	-- ===========================================================================
	function Hz2Time(f_Hz : NATURAL) return TIME is
	begin
		return 1.0 sec / real(f_Hz);
	end function;
	
	function kHz2Time(f_kHz : NATURAL) return TIME is
	begin
		return 1.0 ms / real(f_kHz);
	end function;
	
	function MHz2Time(f_MHz : NATURAL) return TIME
	 is
	begin
		return 1.0 us / real(f_MHz);
	end function;
	
	function GHz2Time(f_GHz : NATURAL) return TIME is
	begin
		return 1.0 ns / real(f_GHz);
	end function;
	
	function THz2Time(f_THz : NATURAL) return TIME is
	begin
		return 1.0 ps / real(f_THz);
	end function;

	
	function Hz2Time(f_Hz : REAL) return TIME is
	begin
		return 1.0 sec / f_Hz;
	end function;
	
	function kHz2Time(f_kHz : REAL) return TIME is
	begin
		return 1.0 ms / f_kHz;
	end function;
	
	function MHz2Time(f_MHz : REAL) return TIME is
	begin
		return 1.0 us / f_MHz;
	end function;
	
	function GHz2Time(f_GHz : REAL) return TIME is
	begin
		return 1.0 ns / f_GHz;
	end function;
	
	function THz2Time(f_THz : REAL) return TIME is
	begin
		return 1.0 ps / f_THz;
	end function;
	
	-- convert standard types (NATURAL, REAL) to frequency (FREQ)
	-- ===========================================================================
	function Hz2Freq(f_Hz : NATURAL) return FREQ is
	begin
		return real(f_Hz) * 1.0 Hz;
	end function;
	
	function kHz2Freq(f_kHz : NATURAL) return FREQ is
	begin
		return real(f_kHz) * 1.0 kHz;
	end function;
	
	function MHz2Freq(f_MHz : NATURAL) return FREQ is
	begin
		return real(f_MHz) * 1.0 MHz;
	end function;
	
	function GHz2Freq(f_GHz : NATURAL) return FREQ is
	begin
		return real(f_GHz) * 1.0 GHz;
	end function;
	
	function THz2Freq(f_THz : NATURAL) return FREQ is
	begin
		return real(f_THz) * 1.0 THz;
	end function;
	
	function Hz2Freq(f_Hz : REAL) return FREQ is
	begin
		return f_Hz * 1.0 Hz;
	end function;
	
	function kHz2Freq(f_kHz : REAL )return FREQ is
	begin
		return f_kHz * 1.0 kHz;
	end function;
	
	function MHz2Freq(f_MHz : REAL )return FREQ is
	begin
		return f_MHz * 1.0 MHz;
	end function;
	
	function GHz2Freq(f_GHz : REAL )return FREQ is
	begin
		return f_GHz * 1.0 GHz;
	end function;
	
	function THz2Freq(f_THz : REAL )return FREQ is
	begin
		return f_THz * 1.0 THz;
	end function;
	
	-- convert TIME to standard type (REAL)
	-- ===========================================================================
	function to_real_fs(t : TIME) return REAL is
	begin
		return real(t / 1.0 fs);
	end;
	
	function to_real_ps(t : TIME) return REAL is
	begin
		return real(t / 1.0 ps);
	end;
	
	function to_real_ns(t : TIME) return REAL is
	begin
		return real(t / 1.0 ns);
	end;
	
	function to_real_us(t : TIME) return REAL is
	begin
		return real(t / 1.0 us);
	end;
	
	function to_real_ms(t : TIME) return REAL is
	begin
		return real(t / 1.0 ms);
	end;
	
	function to_real_sec(t : TIME) return REAL is
	begin
		return real(t / 1.0 sec);
	end;

	-- convert FREQ to standard type (REAL)
	-- ===========================================================================
	function to_real_Hz(f : FREQ) return REAL is
	begin
		return real(f / 1.0 Hz);
	end;
	
	function to_real_kHz(f : FREQ) return REAL is
	begin
		return real(f / 1.0 kHz);
	end;
	
	function to_real_MHz(f : FREQ) return REAL is
	begin
		return real(f / 1.0 MHz);
	end;
	
	function to_real_GHz(f : FREQ) return REAL is
	begin
		return real(f / 1.0 GHz);
	end;
	
	function to_real_THz(f : FREQ) return REAL is
	begin
		return real(f / 1.0 THz);
	end;

	-- convert physical types (TIME, FREQ) to standard type (REAL)
	-- ===========================================================================
	function to_real(t : TIME; scale : TIME) return REAL is
	begin
		if		(scale = 1.0	fs) then	return real(t / 1.0	 fs);
		elsif	(scale = 1.0	ps) then	return real(t / 1.0	 ps);
		elsif	(scale = 1.0	ns) then	return real(t / 1.0	 ns);
		elsif	(scale = 1.0	us) then	return real(t / 1.0	 us);
		elsif	(scale = 1.0	ms) then	return real(t / 1.0	 ms);
		elsif	(scale = 1.0 sec) then	return real(t / 1.0 sec);
		else	report "to_real: scale must have a value of '1.0 <uni>'" severity failure;
		end if;
	end;

	function to_real(f : FREQ; scale : FREQ) return REAL is
	begin
		if		(scale = 1.0	Hz) then	return real(f / 1.0	Hz);
		elsif	(scale = 1.0 kHz) then	return real(f / 1.0 kHz);
		elsif	(scale = 1.0 MHz) then	return real(f / 1.0 MHz);
		elsif	(scale = 1.0 GHz) then	return real(f / 1.0 GHz);
		elsif	(scale = 1.0 THz) then	return real(f / 1.0 THz);
		else	report "to_real: scale must have a value of '1.0 <uni>'" severity failure;
		end if;
	end;

	function to_real(f : BAUD; scale : BAUD) return REAL is
	begin
		if		(scale = 1.0	Bd) then	return real(f / 1.0	 Bd);
		elsif	(scale = 1.0 kBd) then	return real(f / 1.0 kBd);
		elsif	(scale = 1.0 MBd) then	return real(f / 1.0 MBd);
		elsif	(scale = 1.0 GBd) then	return real(f / 1.0 GBd);
		else	report "to_real: scale must have a value of '1.0 <uni>'" severity failure;
		end if;
	end;
	
	function to_real(f : MEMORY; scale : MEMORY) return REAL is
	begin
		if		(scale = 1.0	 B) then	return real(f / 1.0		B);
		elsif	(scale = 1.0 KiB) then	return real(f / 1.0 KiB);
		elsif	(scale = 1.0 MiB) then	return real(f / 1.0 MiB);
		elsif	(scale = 1.0 GiB) then	return real(f / 1.0 GiB);
		elsif	(scale = 1.0 TiB) then	return real(f / 1.0 TiB);
		else	report "to_real: scale must have a value of '1.0 <uni>'" severity failure;
		end if;
	end;
	
	-- calculate needed counter cycles to achieve a given 1. timing/delay and 2. frequency/period
	-- ===========================================================================
	function TimingToCycles(Timing : TIME; Clock_Period : TIME) return NATURAL is
		variable res	: REAL;
	begin
		res := real(Timing / Clock_Period);
		assert not MY_VERBOSE report "TimingToCycles: Timing= " & to_string(Timing) & " Frequency=" & to_string(Clock_Period) & "  return " & str_format(res, 3) severity note;
		return natural(res);
	end;
	
	function TimingToCycles(Timing : TIME; Clock_Frequency : FREQ) return NATURAL is
		variable res	: REAL;
	begin
		res := real(Timing / to_time(Clock_Frequency));
		assert not MY_VERBOSE report "TimingToCycles: Timing= " & to_string(Timing) & " Frequency=" & to_string(Clock_Frequency) & "  return " & str_format(res, 3) severity note;
		return natural(res);
	end;

	-- convert and format physical types to STRING
	function to_string(t : TIME; precision : NATURAL := 3) return STRING is
		variable unit		: STRING(1 to 3)	:= (others => NUL);
		variable value	: REAL;
	begin
		if (t < 1.0 ps) then
			unit(1 to 2)	:= "fs";
			value					:= to_real(t, 1.0 fs);
		elsif (t < 1.0 ns) then
			unit(1 to 2)	:= "ps";
			value					:= to_real(t, 1.0 ps);
		elsif (t < 1.0 us) then
			unit(1 to 2)	:= "ns";
			value					:= to_real(t, 1.0 ns);
		elsif (t < 1.0 ms) then
			unit(1 to 2)	:= "us";
			value					:= to_real(t, 1.0 us);
		elsif (t < 1.0 sec) then
			unit(1 to 2)	:= "ms";
			value					:= to_real(t, 1.0 ms);
		else
			unit					:= "sec";
			value					:= to_real(t, 1.0 sec);
		end if;

		return str_format(value, precision) & " " & str_trim(unit);
	end function;
		
	function to_string(f : FREQ; precision : NATURAL := 3) return STRING is
		variable unit		: STRING(1 to 3)	:= (others => NUL);
		variable value	: REAL;
	begin
		if (f < 1.0 kHz) then
			unit(1 to 2)	:= "Hz";
			value					:= to_real(f, 1.0 Hz);
		elsif (f < 1.0 MHz) then
			unit					:= "kHz";
			value					:= to_real(f, 1.0 kHz);
		elsif (f < 1.0 GHz) then
			unit					:= "MHz";
			value					:= to_real(f, 1.0 MHz);
		elsif (f < 1.0 THz) then
			unit					:= "GHz";
			value					:= to_real(f, 1.0 GHz);
		else
			unit					:= "THz";
			value					:= to_real(f, 1.0 THz);
		end if;

		return str_format(value, precision) & " " & str_trim(unit);
	end function;
		
	function to_string(br : BAUD; precision : NATURAL := 3) return STRING is
		variable unit		: STRING(1 to 3)	:= (others => NUL);
		variable value	: REAL;
	begin
		if (br < 1.0 kBd) then
			unit(1 to 2)	:= "Bd";
			value					:= to_real(br, 1.0 Bd);
		elsif (br < 1.0 MBd) then
			unit					:= "kBd";
			value					:= to_real(br, 1.0 kBd);
		elsif (br < 1.0 GBd) then
			unit					:= "MBd";
			value					:= to_real(br, 1.0 MBd);
		else
			unit					:= "GBd";
			value					:= to_real(br, 1.0 GBd);
		end if;

		return str_format(value, precision) & " " & str_trim(unit);
	end function;
		
	function to_string(mem : MEMORY; precision : NATURAL := 3) return STRING is
		variable unit		: STRING(1 to 3)	:= (others => NUL);
		variable value	: REAL;
	begin
		if (mem < 1.0 KiB) then
			unit(1)				:= 'B';
			value					:= to_real(mem, 1.0 B);
		elsif (mem < 1.0 MiB) then
			unit					:= "KiB";
			value					:= to_real(mem, 1.0 KiB);
		elsif (mem < 1.0 GiB) then
			unit					:= "MiB";
			value					:= to_real(mem, 1.0 MiB);
		elsif (mem < 1.0 TiB) then
			unit					:= "GiB";
			value					:= to_real(mem, 1.0 GiB);
		else
			unit					:= "TiB";
			value					:= to_real(mem, 1.0 TiB);
		end if;

		return str_format(value, precision) & " " & str_trim(unit);
	end function;
	
end package body;
