-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- 
-- ============================================================================
-- Module:				 	TODO
--
-- Authors:				 	Patrick Lehmann
-- 
-- Description:
-- ------------------------------------
--		TODO
--
-- License:
-- ============================================================================
-- Copyright 2007-2014 Technische Universitaet Dresden - Germany
--										 Chair for VLSI-Design, Diagnostics and Architecture
-- 
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
-- 
--		http://www.apache.org/licenses/LICENSE-2.0
-- 
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- ============================================================================


library	IEEE;
use			IEEE.STD_LOGIC_1164.all;

library PoC;
use			PoC.xilinx.all;


entity xil_ChipScopeICON is
	generic (
		PORTS				: POSITIVE
	);
  port (
		ControlBus	: inout	T_CHIPSCOPE_CONTROL_VECTOR(PORTS - 1 downto 0)
	);
end;


architecture rtl of xil_ChipScopeICON is
begin
	assert (PORTS < 16) report "To many ICON control ports." severity failure;

	genICON1 : if (PORTS = 1) generate
		ICON : xil_ChipScopeICON_1
			port map (
				control0		=> ControlBus(0)
			);
	end generate;
	
	genICON2 : if (PORTS = 2) generate
		ICON : xil_ChipScopeICON_2
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1)
			);
	end generate;
	
	genICON3 : if (PORTS = 3) generate
		ICON : xil_ChipScopeICON_3
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2)
			);
	end generate;
	
	genICON4 : if (PORTS = 4) generate
		ICON : xil_ChipScopeICON_4
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3)
			);
	end generate;
	
	genICON5 : if (PORTS = 5) generate
		ICON : xil_ChipScopeICON_5
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4)
			);
	end generate;
	
	genICON6 : if (PORTS = 6) generate
		ICON : xil_ChipScopeICON_6
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4),
				control5		=> ControlBus(5)
			);
	end generate;
	
	genICON7 : if (PORTS = 7) generate
		ICON : xil_ChipScopeICON_7
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4),
				control5		=> ControlBus(5),
				control6		=> ControlBus(6)
			);
	end generate;
	
	genICON8 : if (PORTS = 8) generate
		ICON : xil_ChipScopeICON_8
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4),
				control5		=> ControlBus(5),
				control6		=> ControlBus(6),
				control7		=> ControlBus(7)
			);
	end generate;
	
	genICON9 : if (PORTS = 9) generate
		ICON : xil_ChipScopeICON_9
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4),
				control5		=> ControlBus(5),
				control6		=> ControlBus(6),
				control7		=> ControlBus(7),
				control8		=> ControlBus(8)
			);
	end generate;
	
	genICON10 : if (PORTS = 10) generate
		ICON : xil_ChipScopeICON_10
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4),
				control5		=> ControlBus(5),
				control6		=> ControlBus(6),
				control7		=> ControlBus(7),
				control8		=> ControlBus(8),
				control9		=> ControlBus(9)
			);
	end generate;
	
	genICON11 : if (PORTS = 11) generate
		ICON : xil_ChipScopeICON_11
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4),
				control5		=> ControlBus(5),
				control6		=> ControlBus(6),
				control7		=> ControlBus(7),
				control8		=> ControlBus(8),
				control9		=> ControlBus(9),
				control10		=> ControlBus(10)
			);
	end generate;
	
	genICON12 : if (PORTS = 12) generate
		ICON : xil_ChipScopeICON_12
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4),
				control5		=> ControlBus(5),
				control6		=> ControlBus(6),
				control7		=> ControlBus(7),
				control8		=> ControlBus(8),
				control9		=> ControlBus(9),
				control10		=> ControlBus(10),
				control11		=> ControlBus(11)
			);
	end generate;
	
	genICON13 : if (PORTS = 13) generate
		ICON : xil_ChipScopeICON_13
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4),
				control5		=> ControlBus(5),
				control6		=> ControlBus(6),
				control7		=> ControlBus(7),
				control8		=> ControlBus(8),
				control9		=> ControlBus(9),
				control10		=> ControlBus(10),
				control11		=> ControlBus(11),
				control12		=> ControlBus(12)
			);
	end generate;
	
	genICON14 : if (PORTS = 14) generate
		ICON : xil_ChipScopeICON_14
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4),
				control5		=> ControlBus(5),
				control6		=> ControlBus(6),
				control7		=> ControlBus(7),
				control8		=> ControlBus(8),
				control9		=> ControlBus(9),
				control10		=> ControlBus(10),
				control11		=> ControlBus(11),
				control12		=> ControlBus(12),
				control13		=> ControlBus(13)
			);
	end generate;
	
	genICON15 : if (PORTS = 15) generate
		ICON : xil_ChipScopeICON_15
			port map (
				control0		=> ControlBus(0),
				control1		=> ControlBus(1),
				control2		=> ControlBus(2),
				control3		=> ControlBus(3),
				control4		=> ControlBus(4),
				control5		=> ControlBus(5),
				control6		=> ControlBus(6),
				control7		=> ControlBus(7),
				control8		=> ControlBus(8),
				control9		=> ControlBus(9),
				control10		=> ControlBus(10),
				control11		=> ControlBus(11),
				control12		=> ControlBus(12),
				control13		=> ControlBus(13),
				control14		=> ControlBus(14)
			);
	end generate;
end;
