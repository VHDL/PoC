-- EMACS settings: -*-  tab-width: 2; indent-tabs-mode: t -*-
-- vim: tabstop=2:shiftwidth=2:noexpandtab
-- kate: tab-width 2; replace-tabs off; indent-width 2;
-- =============================================================================
-- Authors:       Gustavo Martin
--
-- Entity:        arith_carrychain_inc_TestHarness
--
-- Description:
-- -------------------------------------
-- Test harness for arith_carrychain_inc component
--
-- License:
-- =============================================================================
-- Copyright 2025-2025 The PoC-Library Authors
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--		http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- =============================================================================

library IEEE;
use     IEEE.std_logic_1164.all;
use     IEEE.numeric_std.all;

library osvvm;
context osvvm.OsvvmContext;

library PoC;


entity arith_carrychain_inc_TestHarness is
end entity;


architecture TestHarness of arith_carrychain_inc_TestHarness is
	constant TPERIOD_CLOCK : time := 10 ns;

	constant BITS : positive := 8;

	signal Clock : std_logic := '1';
	signal Reset : std_logic := '1';

	signal X   : std_logic_vector(BITS - 1 downto 0);
	signal CIn : std_logic;
	signal Y   : std_logic_vector(BITS - 1 downto 0);


	component arith_carrychain_inc_TestController is
		port (
			Clock : in  std_logic;
			Reset : in  std_logic;
			X     : out std_logic_vector;
			CIn   : out std_logic;
			Y     : in  std_logic_vector
		);
	end component;

begin
	Osvvm.ClockResetPkg.CreateClock(
		Clk    => Clock,
		Period => TPERIOD_CLOCK
	);

	Osvvm.ClockResetPkg.CreateReset(
		Reset       => Reset,
		ResetActive => '1',
		Clk         => Clock,
		Period      => 5 * TPERIOD_CLOCK,
		tpd         => 0 ns
	);

	DUT : entity PoC.arith_carrychain_inc
		generic map (
			BITS => BITS
		)
		port map (
			X   => X,
			CIn => CIn,
			Y   => Y
		);

	TestCtrl: component arith_carrychain_inc_TestController
		port map (
			Clock => Clock,
			Reset => Reset,
			X     => X,
			CIn   => CIn,
			Y     => Y
		);

end architecture;
